module mac (CLK,
    rst,
    In1,
    In2,
    MacOut);
 input CLK;
 input rst;
 input [31:0] In1;
 input [31:0] In2;
 output [31:0] MacOut;

 wire \F1.sign_b ;
 wire \In1_reg[0] ;
 wire \In1_reg[10] ;
 wire \In1_reg[11] ;
 wire \In1_reg[12] ;
 wire \In1_reg[13] ;
 wire \In1_reg[14] ;
 wire \In1_reg[15] ;
 wire \In1_reg[16] ;
 wire \In1_reg[17] ;
 wire \In1_reg[18] ;
 wire \In1_reg[19] ;
 wire \In1_reg[1] ;
 wire \In1_reg[20] ;
 wire \In1_reg[21] ;
 wire \In1_reg[22] ;
 wire \In1_reg[2] ;
 wire \In1_reg[31] ;
 wire \In1_reg[3] ;
 wire \In1_reg[4] ;
 wire \In1_reg[5] ;
 wire \In1_reg[6] ;
 wire \In1_reg[7] ;
 wire \In1_reg[8] ;
 wire \In1_reg[9] ;
 wire \In2_reg[0] ;
 wire \In2_reg[10] ;
 wire \In2_reg[12] ;
 wire \In2_reg[14] ;
 wire \In2_reg[16] ;
 wire \In2_reg[18] ;
 wire \In2_reg[20] ;
 wire \In2_reg[22] ;
 wire \In2_reg[2] ;
 wire \In2_reg[31] ;
 wire \In2_reg[4] ;
 wire \In2_reg[6] ;
 wire \In2_reg[8] ;
 wire \M1.U1.U1.u2.instance9_8.Prop_L ;
 wire \M1.U1.U10.u3.instance11_10.Prop_L ;
 wire \M1.U1.U11.u3.instance13_12.Prop_L ;
 wire \M1.U1.U2.u2.instance11_10.Prop_L ;
 wire \M1.U1.U3.u2.instance13_12.Prop_L ;
 wire \M1.U1.U4.u2.instance15_14.Prop_L ;
 wire \M1.U1.U5.u3.instance1_0.Prop_L ;
 wire \M1.U1.U6.u3.instance3_2.Prop_L ;
 wire \M1.U1.U7.u3.instance5_4.Prop_L ;
 wire \M1.U1.U8.u3.instance7_6.Prop_L ;
 wire \M1.U1.U9.u3.instance9_8.Prop_L ;
 wire \M1.ua1.fa0.a ;
 wire \M1.ua1.fa0.b ;
 wire \M1.ua1.fa1.a ;
 wire \M1.ua1.fa1.b ;
 wire \M1.ua1.fa2.a ;
 wire \M1.ua1.fa2.b ;
 wire \M1.ua1.fa3.a ;
 wire \M1.ua1.fa3.b ;
 wire \M1.ua1.fa4.a ;
 wire \M1.ua1.fa4.b ;
 wire \M1.ua1.fa5.a ;
 wire \M1.ua1.fa5.b ;
 wire \M1.ua1.fa6.a ;
 wire \M1.ua1.fa6.b ;
 wire \M1.ua1.fa7.a ;
 wire \M1.ua1.fa7.b ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire clknet_0_CLK;
 wire clknet_3_0__leaf_CLK;
 wire clknet_3_1__leaf_CLK;
 wire clknet_3_2__leaf_CLK;
 wire clknet_3_3__leaf_CLK;
 wire clknet_3_4__leaf_CLK;
 wire clknet_3_5__leaf_CLK;
 wire clknet_3_6__leaf_CLK;
 wire clknet_3_7__leaf_CLK;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;

 sky130_fd_sc_hd__buf_2 _4324_ (.A(net65),
    .X(_1676_));
 sky130_fd_sc_hd__and2_1 _4325_ (.A(_1676_),
    .B(net1),
    .X(_1687_));
 sky130_fd_sc_hd__buf_1 _4326_ (.A(_1687_),
    .X(_0000_));
 sky130_fd_sc_hd__and2_1 _4327_ (.A(_1676_),
    .B(net12),
    .X(_1708_));
 sky130_fd_sc_hd__buf_1 _4328_ (.A(_1708_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_1 _4329_ (.A(_1676_),
    .B(net23),
    .X(_1729_));
 sky130_fd_sc_hd__buf_1 _4330_ (.A(_1729_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _4331_ (.A(_1676_),
    .B(net26),
    .X(_1750_));
 sky130_fd_sc_hd__buf_1 _4332_ (.A(_1750_),
    .X(_0003_));
 sky130_fd_sc_hd__and2_1 _4333_ (.A(_1676_),
    .B(net27),
    .X(_1771_));
 sky130_fd_sc_hd__buf_1 _4334_ (.A(_1771_),
    .X(_0004_));
 sky130_fd_sc_hd__and2_1 _4335_ (.A(_1676_),
    .B(net28),
    .X(_1792_));
 sky130_fd_sc_hd__buf_1 _4336_ (.A(_1792_),
    .X(_0005_));
 sky130_fd_sc_hd__and2_1 _4337_ (.A(_1676_),
    .B(net29),
    .X(_1813_));
 sky130_fd_sc_hd__clkbuf_1 _4338_ (.A(_1813_),
    .X(_0006_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4339_ (.A(net65),
    .X(_1834_));
 sky130_fd_sc_hd__and2_1 _4340_ (.A(_1834_),
    .B(net30),
    .X(_1845_));
 sky130_fd_sc_hd__clkbuf_1 _4341_ (.A(_1845_),
    .X(_0007_));
 sky130_fd_sc_hd__and2_1 _4342_ (.A(_1834_),
    .B(net31),
    .X(_1866_));
 sky130_fd_sc_hd__buf_1 _4343_ (.A(_1866_),
    .X(_0008_));
 sky130_fd_sc_hd__and2_1 _4344_ (.A(_1834_),
    .B(net32),
    .X(_1887_));
 sky130_fd_sc_hd__buf_1 _4345_ (.A(_1887_),
    .X(_0009_));
 sky130_fd_sc_hd__and2_1 _4346_ (.A(_1834_),
    .B(net2),
    .X(_1908_));
 sky130_fd_sc_hd__clkbuf_1 _4347_ (.A(_1908_),
    .X(_0010_));
 sky130_fd_sc_hd__and2_1 _4348_ (.A(_1834_),
    .B(net3),
    .X(_1929_));
 sky130_fd_sc_hd__clkbuf_1 _4349_ (.A(_1929_),
    .X(_0011_));
 sky130_fd_sc_hd__and2_1 _4350_ (.A(_1834_),
    .B(net4),
    .X(_1950_));
 sky130_fd_sc_hd__clkbuf_1 _4351_ (.A(_1950_),
    .X(_0012_));
 sky130_fd_sc_hd__and2_1 _4352_ (.A(_1834_),
    .B(net5),
    .X(_1971_));
 sky130_fd_sc_hd__clkbuf_1 _4353_ (.A(_1971_),
    .X(_0013_));
 sky130_fd_sc_hd__and2_1 _4354_ (.A(_1834_),
    .B(net6),
    .X(_1992_));
 sky130_fd_sc_hd__clkbuf_1 _4355_ (.A(_1992_),
    .X(_0014_));
 sky130_fd_sc_hd__and2_1 _4356_ (.A(_1834_),
    .B(net7),
    .X(_2013_));
 sky130_fd_sc_hd__clkbuf_1 _4357_ (.A(_2013_),
    .X(_0015_));
 sky130_fd_sc_hd__and2_1 _4358_ (.A(_1834_),
    .B(net8),
    .X(_2034_));
 sky130_fd_sc_hd__clkbuf_1 _4359_ (.A(_2034_),
    .X(_0016_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4360_ (.A(net65),
    .X(_2055_));
 sky130_fd_sc_hd__and2_1 _4361_ (.A(_2055_),
    .B(net9),
    .X(_2066_));
 sky130_fd_sc_hd__clkbuf_1 _4362_ (.A(_2066_),
    .X(_0017_));
 sky130_fd_sc_hd__and2_1 _4363_ (.A(_2055_),
    .B(net10),
    .X(_2087_));
 sky130_fd_sc_hd__buf_1 _4364_ (.A(_2087_),
    .X(_0018_));
 sky130_fd_sc_hd__and2_1 _4365_ (.A(_2055_),
    .B(net11),
    .X(_2108_));
 sky130_fd_sc_hd__clkbuf_1 _4366_ (.A(_2108_),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _4367_ (.A(_2055_),
    .B(net13),
    .X(_2129_));
 sky130_fd_sc_hd__buf_1 _4368_ (.A(_2129_),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _4369_ (.A(_2055_),
    .B(net14),
    .X(_2150_));
 sky130_fd_sc_hd__clkbuf_1 _4370_ (.A(_2150_),
    .X(_0021_));
 sky130_fd_sc_hd__and2_1 _4371_ (.A(_2055_),
    .B(net15),
    .X(_2171_));
 sky130_fd_sc_hd__buf_1 _4372_ (.A(_2171_),
    .X(_0022_));
 sky130_fd_sc_hd__and2_1 _4373_ (.A(_2055_),
    .B(net16),
    .X(_2192_));
 sky130_fd_sc_hd__clkbuf_1 _4374_ (.A(_2192_),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _4375_ (.A(_2055_),
    .B(net17),
    .X(_2213_));
 sky130_fd_sc_hd__clkbuf_1 _4376_ (.A(_2213_),
    .X(_0024_));
 sky130_fd_sc_hd__and2_1 _4377_ (.A(_2055_),
    .B(net18),
    .X(_2234_));
 sky130_fd_sc_hd__clkbuf_1 _4378_ (.A(_2234_),
    .X(_0025_));
 sky130_fd_sc_hd__and2_1 _4379_ (.A(_2055_),
    .B(net19),
    .X(_2255_));
 sky130_fd_sc_hd__clkbuf_1 _4380_ (.A(_2255_),
    .X(_0026_));
 sky130_fd_sc_hd__clkbuf_2 _4381_ (.A(net65),
    .X(_2276_));
 sky130_fd_sc_hd__and2_1 _4382_ (.A(_2276_),
    .B(net20),
    .X(_2287_));
 sky130_fd_sc_hd__clkbuf_1 _4383_ (.A(_2287_),
    .X(_0027_));
 sky130_fd_sc_hd__and2_1 _4384_ (.A(_2276_),
    .B(net21),
    .X(_2308_));
 sky130_fd_sc_hd__clkbuf_1 _4385_ (.A(_2308_),
    .X(_0028_));
 sky130_fd_sc_hd__and2_1 _4386_ (.A(_2276_),
    .B(net22),
    .X(_2329_));
 sky130_fd_sc_hd__clkbuf_1 _4387_ (.A(_2329_),
    .X(_0029_));
 sky130_fd_sc_hd__and2_1 _4388_ (.A(_2276_),
    .B(net24),
    .X(_2350_));
 sky130_fd_sc_hd__clkbuf_1 _4389_ (.A(_2350_),
    .X(_0030_));
 sky130_fd_sc_hd__and2_1 _4390_ (.A(_2276_),
    .B(net25),
    .X(_2371_));
 sky130_fd_sc_hd__clkbuf_1 _4391_ (.A(_2371_),
    .X(_0031_));
 sky130_fd_sc_hd__or2_1 _4392_ (.A(\M1.ua1.fa0.b ),
    .B(\M1.ua1.fa0.a ),
    .X(_2392_));
 sky130_fd_sc_hd__nand2_1 _4393_ (.A(\M1.ua1.fa0.b ),
    .B(\M1.ua1.fa0.a ),
    .Y(_2403_));
 sky130_fd_sc_hd__and2_2 _4394_ (.A(_2392_),
    .B(_2403_),
    .X(_2414_));
 sky130_fd_sc_hd__buf_2 _4395_ (.A(\M1.U1.U9.u3.instance9_8.Prop_L ),
    .X(_2425_));
 sky130_fd_sc_hd__buf_2 _4396_ (.A(_2425_),
    .X(_2436_));
 sky130_fd_sc_hd__clkbuf_2 _4397_ (.A(_2436_),
    .X(_2447_));
 sky130_fd_sc_hd__clkbuf_4 _4398_ (.A(_2447_),
    .X(_2458_));
 sky130_fd_sc_hd__clkbuf_4 _4399_ (.A(\In1_reg[21] ),
    .X(_2469_));
 sky130_fd_sc_hd__buf_2 _4400_ (.A(_2469_),
    .X(_2480_));
 sky130_fd_sc_hd__buf_2 _4401_ (.A(_2480_),
    .X(_2491_));
 sky130_fd_sc_hd__nand2_1 _4402_ (.A(_2491_),
    .B(_2458_),
    .Y(_2502_));
 sky130_fd_sc_hd__buf_2 _4403_ (.A(\In2_reg[16] ),
    .X(_2513_));
 sky130_fd_sc_hd__buf_2 _4404_ (.A(_2513_),
    .X(_2524_));
 sky130_fd_sc_hd__clkbuf_2 _4405_ (.A(_2524_),
    .X(_2535_));
 sky130_fd_sc_hd__clkbuf_4 _4406_ (.A(_2535_),
    .X(_2546_));
 sky130_fd_sc_hd__buf_2 _4407_ (.A(\In1_reg[20] ),
    .X(_2557_));
 sky130_fd_sc_hd__buf_2 _4408_ (.A(_2557_),
    .X(_2568_));
 sky130_fd_sc_hd__buf_2 _4409_ (.A(_2568_),
    .X(_2579_));
 sky130_fd_sc_hd__a22o_1 _4410_ (.A1(_2491_),
    .A2(_2546_),
    .B1(_2458_),
    .B2(_2579_),
    .X(_2590_));
 sky130_fd_sc_hd__nand2_1 _4411_ (.A(_2579_),
    .B(_2546_),
    .Y(_2601_));
 sky130_fd_sc_hd__buf_2 _4412_ (.A(\In1_reg[19] ),
    .X(_2612_));
 sky130_fd_sc_hd__buf_2 _4413_ (.A(_2612_),
    .X(_2623_));
 sky130_fd_sc_hd__buf_2 _4414_ (.A(_2623_),
    .X(_2634_));
 sky130_fd_sc_hd__nand2_1 _4415_ (.A(_2634_),
    .B(_2458_),
    .Y(_2645_));
 sky130_fd_sc_hd__xor2_1 _4416_ (.A(_2601_),
    .B(_2645_),
    .X(_2656_));
 sky130_fd_sc_hd__buf_2 _4417_ (.A(\In1_reg[18] ),
    .X(_2667_));
 sky130_fd_sc_hd__buf_2 _4418_ (.A(_2667_),
    .X(_2678_));
 sky130_fd_sc_hd__buf_2 _4419_ (.A(_2678_),
    .X(_2689_));
 sky130_fd_sc_hd__and4_1 _4420_ (.A(_2689_),
    .B(_2634_),
    .C(_2546_),
    .D(_2458_),
    .X(_2700_));
 sky130_fd_sc_hd__buf_2 _4421_ (.A(\In1_reg[17] ),
    .X(_2711_));
 sky130_fd_sc_hd__buf_2 _4422_ (.A(_2711_),
    .X(_2722_));
 sky130_fd_sc_hd__buf_2 _4423_ (.A(_2722_),
    .X(_2733_));
 sky130_fd_sc_hd__and4_1 _4424_ (.A(_2689_),
    .B(_2733_),
    .C(_2535_),
    .D(_2447_),
    .X(_2744_));
 sky130_fd_sc_hd__a22oi_1 _4425_ (.A1(_2689_),
    .A2(_2535_),
    .B1(_2447_),
    .B2(_2733_),
    .Y(_2755_));
 sky130_fd_sc_hd__nor2_1 _4426_ (.A(_2744_),
    .B(_2755_),
    .Y(_2766_));
 sky130_fd_sc_hd__buf_2 _4427_ (.A(\In1_reg[16] ),
    .X(_2777_));
 sky130_fd_sc_hd__buf_2 _4428_ (.A(_2777_),
    .X(_2788_));
 sky130_fd_sc_hd__buf_2 _4429_ (.A(_2788_),
    .X(_2799_));
 sky130_fd_sc_hd__and4_1 _4430_ (.A(_2733_),
    .B(_2799_),
    .C(_2535_),
    .D(_2447_),
    .X(_2810_));
 sky130_fd_sc_hd__buf_2 _4431_ (.A(\In1_reg[15] ),
    .X(_2821_));
 sky130_fd_sc_hd__buf_2 _4432_ (.A(_2821_),
    .X(_2832_));
 sky130_fd_sc_hd__clkbuf_2 _4433_ (.A(_2832_),
    .X(_2843_));
 sky130_fd_sc_hd__buf_2 _4434_ (.A(\In1_reg[14] ),
    .X(_2854_));
 sky130_fd_sc_hd__buf_2 _4435_ (.A(_2854_),
    .X(_2865_));
 sky130_fd_sc_hd__buf_2 _4436_ (.A(_2865_),
    .X(_2876_));
 sky130_fd_sc_hd__a22o_1 _4437_ (.A1(_2843_),
    .A2(_2535_),
    .B1(_2447_),
    .B2(_2876_),
    .X(_2887_));
 sky130_fd_sc_hd__buf_2 _4438_ (.A(\In1_reg[13] ),
    .X(_2898_));
 sky130_fd_sc_hd__buf_2 _4439_ (.A(_2898_),
    .X(_2909_));
 sky130_fd_sc_hd__buf_2 _4440_ (.A(_2909_),
    .X(_2920_));
 sky130_fd_sc_hd__nand2_1 _4441_ (.A(_2920_),
    .B(_2447_),
    .Y(_2931_));
 sky130_fd_sc_hd__nand2_1 _4442_ (.A(_2876_),
    .B(_2535_),
    .Y(_2942_));
 sky130_fd_sc_hd__and4_1 _4443_ (.A(_2876_),
    .B(_2920_),
    .C(_2524_),
    .D(_2436_),
    .X(_2953_));
 sky130_fd_sc_hd__a21o_1 _4444_ (.A1(_2931_),
    .A2(_2942_),
    .B1(_2953_),
    .X(_2964_));
 sky130_fd_sc_hd__clkbuf_2 _4445_ (.A(\In1_reg[12] ),
    .X(_2975_));
 sky130_fd_sc_hd__buf_2 _4446_ (.A(_2975_),
    .X(_2986_));
 sky130_fd_sc_hd__buf_2 _4447_ (.A(_2986_),
    .X(_2997_));
 sky130_fd_sc_hd__a22o_1 _4448_ (.A1(_2920_),
    .A2(_2524_),
    .B1(_2436_),
    .B2(_2997_),
    .X(_3008_));
 sky130_fd_sc_hd__buf_2 _4449_ (.A(\In1_reg[11] ),
    .X(_3019_));
 sky130_fd_sc_hd__buf_2 _4450_ (.A(_3019_),
    .X(_3030_));
 sky130_fd_sc_hd__buf_2 _4451_ (.A(_3030_),
    .X(_3041_));
 sky130_fd_sc_hd__and3_1 _4452_ (.A(_2997_),
    .B(_3041_),
    .C(_2436_),
    .X(_3052_));
 sky130_fd_sc_hd__nand2_1 _4453_ (.A(_3041_),
    .B(_2436_),
    .Y(_3063_));
 sky130_fd_sc_hd__buf_2 _4454_ (.A(\In1_reg[10] ),
    .X(_3074_));
 sky130_fd_sc_hd__buf_2 _4455_ (.A(_3074_),
    .X(_3085_));
 sky130_fd_sc_hd__buf_2 _4456_ (.A(_3085_),
    .X(_3096_));
 sky130_fd_sc_hd__nand2_1 _4457_ (.A(_3096_),
    .B(_2524_),
    .Y(_3107_));
 sky130_fd_sc_hd__buf_2 _4458_ (.A(\In1_reg[9] ),
    .X(_3118_));
 sky130_fd_sc_hd__buf_2 _4459_ (.A(_3118_),
    .X(_3129_));
 sky130_fd_sc_hd__buf_2 _4460_ (.A(_3129_),
    .X(_3140_));
 sky130_fd_sc_hd__and4_1 _4461_ (.A(_3096_),
    .B(_3140_),
    .C(_2524_),
    .D(_2436_),
    .X(_3151_));
 sky130_fd_sc_hd__buf_2 _4462_ (.A(\In1_reg[8] ),
    .X(_3162_));
 sky130_fd_sc_hd__buf_2 _4463_ (.A(_3162_),
    .X(_3173_));
 sky130_fd_sc_hd__buf_2 _4464_ (.A(_3173_),
    .X(_3184_));
 sky130_fd_sc_hd__a22oi_1 _4465_ (.A1(_3140_),
    .A2(_2524_),
    .B1(_2436_),
    .B2(_3184_),
    .Y(_3195_));
 sky130_fd_sc_hd__nand2_1 _4466_ (.A(_3184_),
    .B(_2513_),
    .Y(_3206_));
 sky130_fd_sc_hd__buf_2 _4467_ (.A(\In1_reg[7] ),
    .X(_3217_));
 sky130_fd_sc_hd__buf_2 _4468_ (.A(_3217_),
    .X(_3228_));
 sky130_fd_sc_hd__buf_2 _4469_ (.A(_3228_),
    .X(_3239_));
 sky130_fd_sc_hd__nand2_1 _4470_ (.A(_3239_),
    .B(_2436_),
    .Y(_3250_));
 sky130_fd_sc_hd__and4_1 _4471_ (.A(_3184_),
    .B(_3239_),
    .C(_2513_),
    .D(_2425_),
    .X(_3261_));
 sky130_fd_sc_hd__a21o_1 _4472_ (.A1(_3206_),
    .A2(_3250_),
    .B1(_3261_),
    .X(_3272_));
 sky130_fd_sc_hd__buf_2 _4473_ (.A(\In1_reg[6] ),
    .X(_3283_));
 sky130_fd_sc_hd__buf_2 _4474_ (.A(_3283_),
    .X(_3294_));
 sky130_fd_sc_hd__buf_2 _4475_ (.A(_3294_),
    .X(_3305_));
 sky130_fd_sc_hd__a22o_1 _4476_ (.A1(_3239_),
    .A2(_2513_),
    .B1(_2425_),
    .B2(_3305_),
    .X(_3316_));
 sky130_fd_sc_hd__nand2_1 _4477_ (.A(_3305_),
    .B(_2513_),
    .Y(_3327_));
 sky130_fd_sc_hd__buf_2 _4478_ (.A(\In1_reg[5] ),
    .X(_3338_));
 sky130_fd_sc_hd__buf_2 _4479_ (.A(_3338_),
    .X(_3349_));
 sky130_fd_sc_hd__clkbuf_4 _4480_ (.A(_3349_),
    .X(_3355_));
 sky130_fd_sc_hd__nand2_1 _4481_ (.A(_3355_),
    .B(_2425_),
    .Y(_3362_));
 sky130_fd_sc_hd__and4_1 _4482_ (.A(_3305_),
    .B(_3355_),
    .C(_2513_),
    .D(_2425_),
    .X(_3368_));
 sky130_fd_sc_hd__a21o_1 _4483_ (.A1(_3327_),
    .A2(_3362_),
    .B1(_3368_),
    .X(_3374_));
 sky130_fd_sc_hd__buf_2 _4484_ (.A(\In1_reg[4] ),
    .X(_3380_));
 sky130_fd_sc_hd__buf_2 _4485_ (.A(_3380_),
    .X(_3387_));
 sky130_fd_sc_hd__clkbuf_4 _4486_ (.A(_3387_),
    .X(_3393_));
 sky130_fd_sc_hd__a22o_1 _4487_ (.A1(_3355_),
    .A2(_2513_),
    .B1(_2425_),
    .B2(_3393_),
    .X(_3404_));
 sky130_fd_sc_hd__nand2_1 _4488_ (.A(_3393_),
    .B(_2513_),
    .Y(_3415_));
 sky130_fd_sc_hd__buf_6 _4489_ (.A(\In1_reg[3] ),
    .X(_3426_));
 sky130_fd_sc_hd__buf_2 _4490_ (.A(_3426_),
    .X(_3437_));
 sky130_fd_sc_hd__buf_2 _4491_ (.A(_3437_),
    .X(_3448_));
 sky130_fd_sc_hd__buf_2 _4492_ (.A(_3448_),
    .X(_3459_));
 sky130_fd_sc_hd__nand2_1 _4493_ (.A(_3459_),
    .B(_2425_),
    .Y(_3470_));
 sky130_fd_sc_hd__and4_1 _4494_ (.A(_3393_),
    .B(_3459_),
    .C(\In2_reg[16] ),
    .D(_2425_),
    .X(_3481_));
 sky130_fd_sc_hd__a21oi_1 _4495_ (.A1(_3415_),
    .A2(_3470_),
    .B1(_3481_),
    .Y(_3492_));
 sky130_fd_sc_hd__clkbuf_4 _4496_ (.A(net126),
    .X(_3503_));
 sky130_fd_sc_hd__clkbuf_4 _4497_ (.A(_3503_),
    .X(_3514_));
 sky130_fd_sc_hd__clkbuf_4 _4498_ (.A(_3514_),
    .X(_3525_));
 sky130_fd_sc_hd__buf_6 _4499_ (.A(\In1_reg[0] ),
    .X(_3536_));
 sky130_fd_sc_hd__buf_2 _4500_ (.A(_3536_),
    .X(_3546_));
 sky130_fd_sc_hd__clkbuf_4 _4501_ (.A(_3546_),
    .X(_3556_));
 sky130_fd_sc_hd__and4_1 _4502_ (.A(_3525_),
    .B(_3556_),
    .C(\In2_reg[16] ),
    .D(\M1.U1.U9.u3.instance9_8.Prop_L ),
    .X(_3566_));
 sky130_fd_sc_hd__buf_6 _4503_ (.A(\In1_reg[2] ),
    .X(_3576_));
 sky130_fd_sc_hd__buf_6 _4504_ (.A(_3576_),
    .X(_3586_));
 sky130_fd_sc_hd__buf_2 _4505_ (.A(_3586_),
    .X(_3596_));
 sky130_fd_sc_hd__clkbuf_4 _4506_ (.A(_3596_),
    .X(_3605_));
 sky130_fd_sc_hd__and4_1 _4507_ (.A(_3605_),
    .B(_3525_),
    .C(\In2_reg[16] ),
    .D(\M1.U1.U9.u3.instance9_8.Prop_L ),
    .X(_3616_));
 sky130_fd_sc_hd__and4_1 _4508_ (.A(_3459_),
    .B(_3605_),
    .C(\In2_reg[16] ),
    .D(\M1.U1.U9.u3.instance9_8.Prop_L ),
    .X(_3626_));
 sky130_fd_sc_hd__a211o_1 _4509_ (.A1(_3459_),
    .A2(_3566_),
    .B1(_3616_),
    .C1(_3626_),
    .X(_3635_));
 sky130_fd_sc_hd__a21o_1 _4510_ (.A1(_3492_),
    .A2(_3635_),
    .B1(_3481_),
    .X(_3645_));
 sky130_fd_sc_hd__o2bb2a_1 _4511_ (.A1_N(_3404_),
    .A2_N(_3645_),
    .B1(_3362_),
    .B2(_3415_),
    .X(_3655_));
 sky130_fd_sc_hd__o21bai_1 _4512_ (.A1(_3374_),
    .A2(_3655_),
    .B1_N(_3368_),
    .Y(_3665_));
 sky130_fd_sc_hd__o2bb2a_1 _4513_ (.A1_N(_3316_),
    .A2_N(_3665_),
    .B1(_3250_),
    .B2(_3327_),
    .X(_3675_));
 sky130_fd_sc_hd__o21ba_1 _4514_ (.A1(_3272_),
    .A2(_3675_),
    .B1_N(_3261_),
    .X(_3685_));
 sky130_fd_sc_hd__nand2_1 _4515_ (.A(_3140_),
    .B(_2436_),
    .Y(_3695_));
 sky130_fd_sc_hd__nor2_1 _4516_ (.A(_3695_),
    .B(_3206_),
    .Y(_3704_));
 sky130_fd_sc_hd__o21ba_1 _4517_ (.A1(_3195_),
    .A2(_3685_),
    .B1_N(_3704_),
    .X(_3714_));
 sky130_fd_sc_hd__a21o_1 _4518_ (.A1(_3107_),
    .A2(_3695_),
    .B1(_3151_),
    .X(_3723_));
 sky130_fd_sc_hd__nor2_1 _4519_ (.A(_3714_),
    .B(_3723_),
    .Y(_3732_));
 sky130_fd_sc_hd__or2_1 _4520_ (.A(_3063_),
    .B(_3107_),
    .X(_3742_));
 sky130_fd_sc_hd__a22o_1 _4521_ (.A1(_3041_),
    .A2(_2524_),
    .B1(_2436_),
    .B2(_3096_),
    .X(_3752_));
 sky130_fd_sc_hd__o211a_1 _4522_ (.A1(_3151_),
    .A2(_3732_),
    .B1(_3742_),
    .C1(_3752_),
    .X(_3762_));
 sky130_fd_sc_hd__o21bai_1 _4523_ (.A1(_3063_),
    .A2(_3107_),
    .B1_N(_3762_),
    .Y(_3771_));
 sky130_fd_sc_hd__nand2_1 _4524_ (.A(_2997_),
    .B(_2524_),
    .Y(_3781_));
 sky130_fd_sc_hd__nand2_1 _4525_ (.A(_3781_),
    .B(_3063_),
    .Y(_3783_));
 sky130_fd_sc_hd__a22o_1 _4526_ (.A1(_2524_),
    .A2(_3052_),
    .B1(_3771_),
    .B2(_3783_),
    .X(_3784_));
 sky130_fd_sc_hd__o2bb2a_1 _4527_ (.A1_N(_3008_),
    .A2_N(_3784_),
    .B1(_2931_),
    .B2(_3781_),
    .X(_3785_));
 sky130_fd_sc_hd__nor2_1 _4528_ (.A(_2964_),
    .B(_3785_),
    .Y(_3786_));
 sky130_fd_sc_hd__and4_1 _4529_ (.A(_2843_),
    .B(_2876_),
    .C(_2535_),
    .D(_2447_),
    .X(_3787_));
 sky130_fd_sc_hd__a211o_1 _4530_ (.A1(_2887_),
    .A2(_3786_),
    .B1(_3787_),
    .C1(_2953_),
    .X(_3788_));
 sky130_fd_sc_hd__a22o_1 _4531_ (.A1(_2799_),
    .A2(_2535_),
    .B1(_2447_),
    .B2(_2843_),
    .X(_3789_));
 sky130_fd_sc_hd__and4_1 _4532_ (.A(_2799_),
    .B(_2843_),
    .C(_2535_),
    .D(_2447_),
    .X(_3790_));
 sky130_fd_sc_hd__a21o_1 _4533_ (.A1(_3788_),
    .A2(_3789_),
    .B1(_3790_),
    .X(_3791_));
 sky130_fd_sc_hd__a22o_1 _4534_ (.A1(_2733_),
    .A2(_2535_),
    .B1(_2447_),
    .B2(_2799_),
    .X(_3792_));
 sky130_fd_sc_hd__o21a_1 _4535_ (.A1(_2810_),
    .A2(_3791_),
    .B1(_3792_),
    .X(_3793_));
 sky130_fd_sc_hd__a21o_1 _4536_ (.A1(_2766_),
    .A2(_3793_),
    .B1(_2744_),
    .X(_3794_));
 sky130_fd_sc_hd__a22o_1 _4537_ (.A1(_2634_),
    .A2(_2546_),
    .B1(_2458_),
    .B2(_2689_),
    .X(_3795_));
 sky130_fd_sc_hd__o21a_1 _4538_ (.A1(_2700_),
    .A2(_3794_),
    .B1(_3795_),
    .X(_3796_));
 sky130_fd_sc_hd__a2bb2oi_1 _4539_ (.A1_N(_2601_),
    .A2_N(_2645_),
    .B1(_2656_),
    .B2(_3796_),
    .Y(_3797_));
 sky130_fd_sc_hd__inv_2 _4540_ (.A(_3797_),
    .Y(_3798_));
 sky130_fd_sc_hd__o2bb2a_1 _4541_ (.A1_N(_2590_),
    .A2_N(_3798_),
    .B1(_2502_),
    .B2(_2601_),
    .X(_3799_));
 sky130_fd_sc_hd__buf_2 _4542_ (.A(\In1_reg[22] ),
    .X(_3800_));
 sky130_fd_sc_hd__buf_2 _4543_ (.A(_3800_),
    .X(_3801_));
 sky130_fd_sc_hd__and3_1 _4544_ (.A(_3801_),
    .B(_2546_),
    .C(_2458_),
    .X(_3802_));
 sky130_fd_sc_hd__o21ba_1 _4545_ (.A1(_2502_),
    .A2(_3799_),
    .B1_N(_3802_),
    .X(_3803_));
 sky130_fd_sc_hd__buf_2 _4546_ (.A(_2579_),
    .X(_3804_));
 sky130_fd_sc_hd__buf_2 _4547_ (.A(\M1.U1.U10.u3.instance11_10.Prop_L ),
    .X(_3805_));
 sky130_fd_sc_hd__buf_2 _4548_ (.A(_3805_),
    .X(_3806_));
 sky130_fd_sc_hd__clkbuf_2 _4549_ (.A(_3806_),
    .X(_3807_));
 sky130_fd_sc_hd__buf_2 _4550_ (.A(_3807_),
    .X(_3808_));
 sky130_fd_sc_hd__buf_2 _4551_ (.A(\In2_reg[18] ),
    .X(_3809_));
 sky130_fd_sc_hd__buf_2 _4552_ (.A(_3809_),
    .X(_3810_));
 sky130_fd_sc_hd__clkbuf_2 _4553_ (.A(_3810_),
    .X(_3811_));
 sky130_fd_sc_hd__buf_2 _4554_ (.A(_3811_),
    .X(_3812_));
 sky130_fd_sc_hd__a22o_1 _4555_ (.A1(_3804_),
    .A2(_3808_),
    .B1(_3812_),
    .B2(_2491_),
    .X(_3813_));
 sky130_fd_sc_hd__buf_2 _4556_ (.A(_2634_),
    .X(_3814_));
 sky130_fd_sc_hd__nand2_1 _4557_ (.A(_3814_),
    .B(_3808_),
    .Y(_3815_));
 sky130_fd_sc_hd__nand2_1 _4558_ (.A(_3804_),
    .B(_3812_),
    .Y(_3816_));
 sky130_fd_sc_hd__and4_1 _4559_ (.A(_3804_),
    .B(_3814_),
    .C(_3808_),
    .D(_3812_),
    .X(_3817_));
 sky130_fd_sc_hd__a21o_1 _4560_ (.A1(_3815_),
    .A2(_3816_),
    .B1(_3817_),
    .X(_3818_));
 sky130_fd_sc_hd__buf_2 _4561_ (.A(_2689_),
    .X(_3819_));
 sky130_fd_sc_hd__a22o_1 _4562_ (.A1(_3819_),
    .A2(_3808_),
    .B1(_3812_),
    .B2(_3814_),
    .X(_3820_));
 sky130_fd_sc_hd__nand2_1 _4563_ (.A(_3819_),
    .B(_3812_),
    .Y(_3821_));
 sky130_fd_sc_hd__clkbuf_2 _4564_ (.A(_2733_),
    .X(_3822_));
 sky130_fd_sc_hd__nand2_1 _4565_ (.A(_3822_),
    .B(_3808_),
    .Y(_3823_));
 sky130_fd_sc_hd__and4_1 _4566_ (.A(_3819_),
    .B(_3822_),
    .C(_3807_),
    .D(_3812_),
    .X(_3824_));
 sky130_fd_sc_hd__a21o_1 _4567_ (.A1(_3821_),
    .A2(_3823_),
    .B1(_3824_),
    .X(_3825_));
 sky130_fd_sc_hd__clkbuf_2 _4568_ (.A(_2799_),
    .X(_3826_));
 sky130_fd_sc_hd__and4_1 _4569_ (.A(_2733_),
    .B(_3826_),
    .C(_3807_),
    .D(_3811_),
    .X(_3827_));
 sky130_fd_sc_hd__clkbuf_2 _4570_ (.A(_2843_),
    .X(_3828_));
 sky130_fd_sc_hd__and4_1 _4571_ (.A(_2799_),
    .B(_3828_),
    .C(_3807_),
    .D(_3811_),
    .X(_3829_));
 sky130_fd_sc_hd__a22oi_1 _4572_ (.A1(_3828_),
    .A2(_3807_),
    .B1(_3811_),
    .B2(_3826_),
    .Y(_3830_));
 sky130_fd_sc_hd__nor2_1 _4573_ (.A(_3829_),
    .B(_3830_),
    .Y(_3831_));
 sky130_fd_sc_hd__clkbuf_2 _4574_ (.A(_2876_),
    .X(_3832_));
 sky130_fd_sc_hd__and4_1 _4575_ (.A(_2843_),
    .B(_3832_),
    .C(_3807_),
    .D(_3811_),
    .X(_3833_));
 sky130_fd_sc_hd__buf_2 _4576_ (.A(_3041_),
    .X(_3834_));
 sky130_fd_sc_hd__and4_1 _4577_ (.A(_2997_),
    .B(_3834_),
    .C(_3806_),
    .D(_3810_),
    .X(_3835_));
 sky130_fd_sc_hd__buf_2 _4578_ (.A(_2997_),
    .X(_3836_));
 sky130_fd_sc_hd__a22oi_1 _4579_ (.A1(_3834_),
    .A2(_3806_),
    .B1(_3810_),
    .B2(_3836_),
    .Y(_3837_));
 sky130_fd_sc_hd__or2_1 _4580_ (.A(_3835_),
    .B(_3837_),
    .X(_3838_));
 sky130_fd_sc_hd__and4_1 _4581_ (.A(_2920_),
    .B(_3836_),
    .C(_3806_),
    .D(_3810_),
    .X(_3839_));
 sky130_fd_sc_hd__clkbuf_2 _4582_ (.A(_2920_),
    .X(_3840_));
 sky130_fd_sc_hd__a22oi_1 _4583_ (.A1(_3836_),
    .A2(_3806_),
    .B1(_3811_),
    .B2(_3840_),
    .Y(_3841_));
 sky130_fd_sc_hd__or2_1 _4584_ (.A(_3839_),
    .B(_3841_),
    .X(_3842_));
 sky130_fd_sc_hd__nor2_1 _4585_ (.A(_3838_),
    .B(_3842_),
    .Y(_3843_));
 sky130_fd_sc_hd__buf_2 _4586_ (.A(_3096_),
    .X(_3844_));
 sky130_fd_sc_hd__and4_1 _4587_ (.A(_3041_),
    .B(_3844_),
    .C(_3806_),
    .D(_3810_),
    .X(_3845_));
 sky130_fd_sc_hd__a22oi_1 _4588_ (.A1(_3844_),
    .A2(_3806_),
    .B1(_3810_),
    .B2(_3834_),
    .Y(_3846_));
 sky130_fd_sc_hd__or2_1 _4589_ (.A(_3845_),
    .B(_3846_),
    .X(_3847_));
 sky130_fd_sc_hd__buf_2 _4590_ (.A(_3184_),
    .X(_3848_));
 sky130_fd_sc_hd__buf_2 _4591_ (.A(_3140_),
    .X(_3849_));
 sky130_fd_sc_hd__a22o_1 _4592_ (.A1(_3848_),
    .A2(_3806_),
    .B1(_3810_),
    .B2(_3849_),
    .X(_3850_));
 sky130_fd_sc_hd__buf_2 _4593_ (.A(_3239_),
    .X(_3851_));
 sky130_fd_sc_hd__nand2_1 _4594_ (.A(_3851_),
    .B(_3805_),
    .Y(_3852_));
 sky130_fd_sc_hd__buf_2 _4595_ (.A(_3305_),
    .X(_3853_));
 sky130_fd_sc_hd__nand2_1 _4596_ (.A(_3853_),
    .B(_3809_),
    .Y(_3854_));
 sky130_fd_sc_hd__a22o_1 _4597_ (.A1(_3853_),
    .A2(_3805_),
    .B1(_3809_),
    .B2(_3851_),
    .X(_3855_));
 sky130_fd_sc_hd__o21a_1 _4598_ (.A1(_3852_),
    .A2(_3854_),
    .B1(_3855_),
    .X(_3856_));
 sky130_fd_sc_hd__clkbuf_2 _4599_ (.A(_3355_),
    .X(_3857_));
 sky130_fd_sc_hd__and4_1 _4600_ (.A(_3853_),
    .B(_3857_),
    .C(_3805_),
    .D(_3809_),
    .X(_3858_));
 sky130_fd_sc_hd__clkbuf_2 _4601_ (.A(_3393_),
    .X(_3859_));
 sky130_fd_sc_hd__a22o_1 _4602_ (.A1(_3859_),
    .A2(_3805_),
    .B1(_3809_),
    .B2(_3355_),
    .X(_3860_));
 sky130_fd_sc_hd__nand2_1 _4603_ (.A(_3859_),
    .B(_3809_),
    .Y(_3861_));
 sky130_fd_sc_hd__clkbuf_2 _4604_ (.A(_3459_),
    .X(_3862_));
 sky130_fd_sc_hd__nand2_1 _4605_ (.A(_3862_),
    .B(\M1.U1.U10.u3.instance11_10.Prop_L ),
    .Y(_3863_));
 sky130_fd_sc_hd__and4_1 _4606_ (.A(_3393_),
    .B(_3459_),
    .C(\M1.U1.U10.u3.instance11_10.Prop_L ),
    .D(_3809_),
    .X(_3864_));
 sky130_fd_sc_hd__a21o_1 _4607_ (.A1(_3861_),
    .A2(_3863_),
    .B1(_3864_),
    .X(_3865_));
 sky130_fd_sc_hd__a22o_1 _4608_ (.A1(_3605_),
    .A2(\M1.U1.U10.u3.instance11_10.Prop_L ),
    .B1(_3809_),
    .B2(_3459_),
    .X(_3866_));
 sky130_fd_sc_hd__inv_2 _4609_ (.A(_3525_),
    .Y(_3867_));
 sky130_fd_sc_hd__nand2_1 _4610_ (.A(_3605_),
    .B(\In2_reg[18] ),
    .Y(_3868_));
 sky130_fd_sc_hd__nor2_1 _4611_ (.A(_3867_),
    .B(_3868_),
    .Y(_3869_));
 sky130_fd_sc_hd__nand2_1 _4612_ (.A(_3525_),
    .B(\M1.U1.U10.u3.instance11_10.Prop_L ),
    .Y(_3870_));
 sky130_fd_sc_hd__nand2_1 _4613_ (.A(_3556_),
    .B(\In2_reg[18] ),
    .Y(_3871_));
 sky130_fd_sc_hd__or2_1 _4614_ (.A(_3870_),
    .B(_3871_),
    .X(_3872_));
 sky130_fd_sc_hd__a21bo_1 _4615_ (.A1(\M1.U1.U10.u3.instance11_10.Prop_L ),
    .A2(_3869_),
    .B1_N(_3872_),
    .X(_3873_));
 sky130_fd_sc_hd__o2bb2a_1 _4616_ (.A1_N(_3866_),
    .A2_N(_3873_),
    .B1(_3863_),
    .B2(_3868_),
    .X(_3874_));
 sky130_fd_sc_hd__o21bai_1 _4617_ (.A1(_3865_),
    .A2(_3874_),
    .B1_N(_3864_),
    .Y(_3875_));
 sky130_fd_sc_hd__nand2_1 _4618_ (.A(_3857_),
    .B(_3805_),
    .Y(_3876_));
 sky130_fd_sc_hd__o2bb2a_1 _4619_ (.A1_N(_3860_),
    .A2_N(_3875_),
    .B1(_3876_),
    .B2(_3861_),
    .X(_3877_));
 sky130_fd_sc_hd__a21o_1 _4620_ (.A1(_3854_),
    .A2(_3876_),
    .B1(_3858_),
    .X(_3878_));
 sky130_fd_sc_hd__nor2_1 _4621_ (.A(_3877_),
    .B(_3878_),
    .Y(_3879_));
 sky130_fd_sc_hd__or2_1 _4622_ (.A(_3858_),
    .B(_3879_),
    .X(_3880_));
 sky130_fd_sc_hd__nor2_1 _4623_ (.A(_3852_),
    .B(_3854_),
    .Y(_3881_));
 sky130_fd_sc_hd__a21oi_1 _4624_ (.A1(_3856_),
    .A2(_3880_),
    .B1(_3881_),
    .Y(_3882_));
 sky130_fd_sc_hd__and3_1 _4625_ (.A(_3848_),
    .B(_3851_),
    .C(_3809_),
    .X(_3883_));
 sky130_fd_sc_hd__nand2_1 _4626_ (.A(_3848_),
    .B(_3810_),
    .Y(_3884_));
 sky130_fd_sc_hd__a22o_1 _4627_ (.A1(_3805_),
    .A2(_3883_),
    .B1(_3852_),
    .B2(_3884_),
    .X(_3885_));
 sky130_fd_sc_hd__a2bb2o_1 _4628_ (.A1_N(_3882_),
    .A2_N(_3885_),
    .B1(_3805_),
    .B2(_3883_),
    .X(_3886_));
 sky130_fd_sc_hd__nand2_1 _4629_ (.A(_3849_),
    .B(_3806_),
    .Y(_3887_));
 sky130_fd_sc_hd__o2bb2a_1 _4630_ (.A1_N(_3850_),
    .A2_N(_3886_),
    .B1(_3884_),
    .B2(_3887_),
    .X(_3888_));
 sky130_fd_sc_hd__nand2_1 _4631_ (.A(_3844_),
    .B(_3810_),
    .Y(_3889_));
 sky130_fd_sc_hd__and4_1 _4632_ (.A(_3096_),
    .B(_3849_),
    .C(_3806_),
    .D(_3810_),
    .X(_3890_));
 sky130_fd_sc_hd__a21o_1 _4633_ (.A1(_3889_),
    .A2(_3887_),
    .B1(_3890_),
    .X(_3891_));
 sky130_fd_sc_hd__o21ba_1 _4634_ (.A1(_3888_),
    .A2(_3891_),
    .B1_N(_3890_),
    .X(_3892_));
 sky130_fd_sc_hd__o21ba_1 _4635_ (.A1(_3847_),
    .A2(_3892_),
    .B1_N(_3845_),
    .X(_3893_));
 sky130_fd_sc_hd__inv_2 _4636_ (.A(_3893_),
    .Y(_3894_));
 sky130_fd_sc_hd__a211oi_1 _4637_ (.A1(_3843_),
    .A2(_3894_),
    .B1(_3835_),
    .C1(_3839_),
    .Y(_3895_));
 sky130_fd_sc_hd__a22oi_1 _4638_ (.A1(_3840_),
    .A2(_3807_),
    .B1(_3811_),
    .B2(_3832_),
    .Y(_3896_));
 sky130_fd_sc_hd__and4_1 _4639_ (.A(_2876_),
    .B(_3840_),
    .C(_3807_),
    .D(_3811_),
    .X(_3897_));
 sky130_fd_sc_hd__o21bai_1 _4640_ (.A1(_3895_),
    .A2(_3896_),
    .B1_N(_3897_),
    .Y(_3898_));
 sky130_fd_sc_hd__a22o_1 _4641_ (.A1(_3832_),
    .A2(_3807_),
    .B1(_3811_),
    .B2(_3828_),
    .X(_3899_));
 sky130_fd_sc_hd__o21a_1 _4642_ (.A1(_3833_),
    .A2(_3898_),
    .B1(_3899_),
    .X(_3900_));
 sky130_fd_sc_hd__a21o_1 _4643_ (.A1(_3831_),
    .A2(_3900_),
    .B1(_3829_),
    .X(_3901_));
 sky130_fd_sc_hd__a22o_1 _4644_ (.A1(_3826_),
    .A2(_3807_),
    .B1(_3811_),
    .B2(_3822_),
    .X(_3902_));
 sky130_fd_sc_hd__o21ai_1 _4645_ (.A1(_3827_),
    .A2(_3901_),
    .B1(_3902_),
    .Y(_3903_));
 sky130_fd_sc_hd__o21bai_1 _4646_ (.A1(_3825_),
    .A2(_3903_),
    .B1_N(_3824_),
    .Y(_3904_));
 sky130_fd_sc_hd__o2bb2a_1 _4647_ (.A1_N(_3820_),
    .A2_N(_3904_),
    .B1(_3815_),
    .B2(_3821_),
    .X(_3905_));
 sky130_fd_sc_hd__nor2_1 _4648_ (.A(_3818_),
    .B(_3905_),
    .Y(_3906_));
 sky130_fd_sc_hd__buf_2 _4649_ (.A(_2491_),
    .X(_3907_));
 sky130_fd_sc_hd__nand2_1 _4650_ (.A(_3907_),
    .B(_3808_),
    .Y(_3908_));
 sky130_fd_sc_hd__nor2_1 _4651_ (.A(_3816_),
    .B(_3908_),
    .Y(_3909_));
 sky130_fd_sc_hd__a211o_1 _4652_ (.A1(_3813_),
    .A2(_3906_),
    .B1(_3909_),
    .C1(_3817_),
    .X(_3910_));
 sky130_fd_sc_hd__buf_2 _4653_ (.A(_3801_),
    .X(_3911_));
 sky130_fd_sc_hd__a21boi_1 _4654_ (.A1(_3911_),
    .A2(_3812_),
    .B1_N(_3908_),
    .Y(_3912_));
 sky130_fd_sc_hd__and4_1 _4655_ (.A(_3911_),
    .B(_3907_),
    .C(_3808_),
    .D(_3812_),
    .X(_3913_));
 sky130_fd_sc_hd__nor2_1 _4656_ (.A(_3912_),
    .B(_3913_),
    .Y(_3914_));
 sky130_fd_sc_hd__and2_1 _4657_ (.A(_3910_),
    .B(_3914_),
    .X(_3915_));
 sky130_fd_sc_hd__nor2_1 _4658_ (.A(_3910_),
    .B(_3914_),
    .Y(_3916_));
 sky130_fd_sc_hd__nor2_1 _4659_ (.A(_3915_),
    .B(_3916_),
    .Y(_3917_));
 sky130_fd_sc_hd__and3_1 _4660_ (.A(_2458_),
    .B(_3803_),
    .C(_3917_),
    .X(_3918_));
 sky130_fd_sc_hd__o21ai_1 _4661_ (.A1(_3816_),
    .A2(_3908_),
    .B1(_3813_),
    .Y(_3919_));
 sky130_fd_sc_hd__or2_1 _4662_ (.A(_3817_),
    .B(_3906_),
    .X(_3920_));
 sky130_fd_sc_hd__xnor2_1 _4663_ (.A(_3919_),
    .B(_3920_),
    .Y(_3921_));
 sky130_fd_sc_hd__a21boi_1 _4664_ (.A1(_3911_),
    .A2(_2546_),
    .B1_N(_2502_),
    .Y(_3922_));
 sky130_fd_sc_hd__a21oi_1 _4665_ (.A1(_2491_),
    .A2(_3802_),
    .B1(_3922_),
    .Y(_3923_));
 sky130_fd_sc_hd__nor2b_1 _4666_ (.A(_3799_),
    .B_N(_3923_),
    .Y(_3924_));
 sky130_fd_sc_hd__a21oi_1 _4667_ (.A1(_3911_),
    .A2(_2458_),
    .B1(_2546_),
    .Y(_3925_));
 sky130_fd_sc_hd__a21o_1 _4668_ (.A1(_3907_),
    .A2(_3802_),
    .B1(_3924_),
    .X(_3926_));
 sky130_fd_sc_hd__o21ai_1 _4669_ (.A1(_3802_),
    .A2(_3925_),
    .B1(_3926_),
    .Y(_3927_));
 sky130_fd_sc_hd__o31ai_1 _4670_ (.A1(_3802_),
    .A2(_3924_),
    .A3(_3925_),
    .B1(_3927_),
    .Y(_3928_));
 sky130_fd_sc_hd__nand2_1 _4671_ (.A(_3921_),
    .B(_3928_),
    .Y(_3929_));
 sky130_fd_sc_hd__and2b_1 _4672_ (.A_N(_3923_),
    .B(_3799_),
    .X(_3930_));
 sky130_fd_sc_hd__nor2_1 _4673_ (.A(_3924_),
    .B(_3930_),
    .Y(_3931_));
 sky130_fd_sc_hd__inv_2 _4674_ (.A(_3931_),
    .Y(_3932_));
 sky130_fd_sc_hd__and2_1 _4675_ (.A(_3818_),
    .B(_3905_),
    .X(_3933_));
 sky130_fd_sc_hd__or2_1 _4676_ (.A(_3906_),
    .B(_3933_),
    .X(_3934_));
 sky130_fd_sc_hd__nor2_1 _4677_ (.A(_3932_),
    .B(_3934_),
    .Y(_3935_));
 sky130_fd_sc_hd__and2_1 _4678_ (.A(_3932_),
    .B(_3934_),
    .X(_3936_));
 sky130_fd_sc_hd__or2_1 _4679_ (.A(_3935_),
    .B(_3936_),
    .X(_3937_));
 sky130_fd_sc_hd__o21a_1 _4680_ (.A1(_2502_),
    .A2(_2601_),
    .B1(_2590_),
    .X(_3938_));
 sky130_fd_sc_hd__xnor2_1 _4681_ (.A(_3938_),
    .B(_3797_),
    .Y(_3939_));
 sky130_fd_sc_hd__inv_2 _4682_ (.A(_3939_),
    .Y(_3940_));
 sky130_fd_sc_hd__o21a_1 _4683_ (.A1(_3815_),
    .A2(_3821_),
    .B1(_3820_),
    .X(_3941_));
 sky130_fd_sc_hd__xnor2_1 _4684_ (.A(_3941_),
    .B(_3904_),
    .Y(_3942_));
 sky130_fd_sc_hd__nor2_1 _4685_ (.A(_3940_),
    .B(_3942_),
    .Y(_3943_));
 sky130_fd_sc_hd__and2_1 _4686_ (.A(_3940_),
    .B(_3942_),
    .X(_3944_));
 sky130_fd_sc_hd__or2_1 _4687_ (.A(_3943_),
    .B(_3944_),
    .X(_3945_));
 sky130_fd_sc_hd__xnor2_1 _4688_ (.A(_2656_),
    .B(_3796_),
    .Y(_3946_));
 sky130_fd_sc_hd__xnor2_1 _4689_ (.A(_3825_),
    .B(_3903_),
    .Y(_3947_));
 sky130_fd_sc_hd__inv_2 _4690_ (.A(_3795_),
    .Y(_3948_));
 sky130_fd_sc_hd__nor2_1 _4691_ (.A(_3948_),
    .B(_2700_),
    .Y(_3949_));
 sky130_fd_sc_hd__xor2_1 _4692_ (.A(_3794_),
    .B(_3949_),
    .X(_3950_));
 sky130_fd_sc_hd__or2b_1 _4693_ (.A(_3827_),
    .B_N(_3902_),
    .X(_3951_));
 sky130_fd_sc_hd__xnor2_1 _4694_ (.A(_3901_),
    .B(_3951_),
    .Y(_3952_));
 sky130_fd_sc_hd__and2_1 _4695_ (.A(_3950_),
    .B(_3952_),
    .X(_3953_));
 sky130_fd_sc_hd__xor2_1 _4696_ (.A(_2766_),
    .B(_3793_),
    .X(_3954_));
 sky130_fd_sc_hd__xor2_1 _4697_ (.A(_3831_),
    .B(_3900_),
    .X(_3955_));
 sky130_fd_sc_hd__and2_1 _4698_ (.A(_3954_),
    .B(_3955_),
    .X(_3956_));
 sky130_fd_sc_hd__inv_2 _4699_ (.A(_2810_),
    .Y(_3957_));
 sky130_fd_sc_hd__nand2_1 _4700_ (.A(_3792_),
    .B(_3957_),
    .Y(_3958_));
 sky130_fd_sc_hd__xnor2_1 _4701_ (.A(_3791_),
    .B(_3958_),
    .Y(_3959_));
 sky130_fd_sc_hd__nand2_1 _4702_ (.A(_3833_),
    .B(_3898_),
    .Y(_3960_));
 sky130_fd_sc_hd__o2bb2a_1 _4703_ (.A1_N(_3900_),
    .A2_N(_3960_),
    .B1(_3899_),
    .B2(_3898_),
    .X(_3961_));
 sky130_fd_sc_hd__nand2_1 _4704_ (.A(_3959_),
    .B(_3961_),
    .Y(_3962_));
 sky130_fd_sc_hd__and2b_1 _4705_ (.A_N(_3790_),
    .B(_3789_),
    .X(_3963_));
 sky130_fd_sc_hd__xnor2_1 _4706_ (.A(_3788_),
    .B(_3963_),
    .Y(_3964_));
 sky130_fd_sc_hd__nor2_1 _4707_ (.A(_3897_),
    .B(_3896_),
    .Y(_3965_));
 sky130_fd_sc_hd__xnor2_1 _4708_ (.A(_3895_),
    .B(_3965_),
    .Y(_3966_));
 sky130_fd_sc_hd__and2b_1 _4709_ (.A_N(_3964_),
    .B(_3966_),
    .X(_3967_));
 sky130_fd_sc_hd__inv_2 _4710_ (.A(_3787_),
    .Y(_3968_));
 sky130_fd_sc_hd__a211o_1 _4711_ (.A1(_2887_),
    .A2(_3968_),
    .B1(_3786_),
    .C1(_2953_),
    .X(_3969_));
 sky130_fd_sc_hd__o211ai_1 _4712_ (.A1(_2953_),
    .A2(_3786_),
    .B1(_3968_),
    .C1(_2887_),
    .Y(_3970_));
 sky130_fd_sc_hd__nand2_1 _4713_ (.A(_3969_),
    .B(_3970_),
    .Y(_3971_));
 sky130_fd_sc_hd__o21ba_1 _4714_ (.A1(_3838_),
    .A2(_3893_),
    .B1_N(_3835_),
    .X(_3972_));
 sky130_fd_sc_hd__xnor2_1 _4715_ (.A(_3842_),
    .B(_3972_),
    .Y(_3973_));
 sky130_fd_sc_hd__nor2_1 _4716_ (.A(_3971_),
    .B(_3973_),
    .Y(_3974_));
 sky130_fd_sc_hd__and2_1 _4717_ (.A(_2964_),
    .B(_3785_),
    .X(_3975_));
 sky130_fd_sc_hd__or2_1 _4718_ (.A(_3786_),
    .B(_3975_),
    .X(_3976_));
 sky130_fd_sc_hd__xnor2_1 _4719_ (.A(_3838_),
    .B(_3893_),
    .Y(_3977_));
 sky130_fd_sc_hd__or2_1 _4720_ (.A(_3976_),
    .B(_3977_),
    .X(_3978_));
 sky130_fd_sc_hd__o21a_1 _4721_ (.A1(_2931_),
    .A2(_3781_),
    .B1(_3008_),
    .X(_3979_));
 sky130_fd_sc_hd__xnor2_1 _4722_ (.A(_3979_),
    .B(_3784_),
    .Y(_3980_));
 sky130_fd_sc_hd__xnor2_1 _4723_ (.A(_3847_),
    .B(_3892_),
    .Y(_3981_));
 sky130_fd_sc_hd__nor2_1 _4724_ (.A(_3980_),
    .B(_3981_),
    .Y(_3982_));
 sky130_fd_sc_hd__a22o_1 _4725_ (.A1(_3781_),
    .A2(_3063_),
    .B1(_3052_),
    .B2(_2524_),
    .X(_3983_));
 sky130_fd_sc_hd__xnor2_1 _4726_ (.A(_3771_),
    .B(_3983_),
    .Y(_3984_));
 sky130_fd_sc_hd__xor2_1 _4727_ (.A(_3888_),
    .B(_3891_),
    .X(_3985_));
 sky130_fd_sc_hd__and2_1 _4728_ (.A(_3984_),
    .B(_3985_),
    .X(_3986_));
 sky130_fd_sc_hd__a211oi_1 _4729_ (.A1(_3742_),
    .A2(_3752_),
    .B1(_3151_),
    .C1(_3732_),
    .Y(_3987_));
 sky130_fd_sc_hd__or2_1 _4730_ (.A(_3762_),
    .B(_3987_),
    .X(_3988_));
 sky130_fd_sc_hd__o21a_1 _4731_ (.A1(_3884_),
    .A2(_3887_),
    .B1(_3850_),
    .X(_3989_));
 sky130_fd_sc_hd__xnor2_1 _4732_ (.A(_3989_),
    .B(_3886_),
    .Y(_3990_));
 sky130_fd_sc_hd__or2_1 _4733_ (.A(_3988_),
    .B(_3990_),
    .X(_3991_));
 sky130_fd_sc_hd__xor2_1 _4734_ (.A(_3714_),
    .B(_3723_),
    .X(_3992_));
 sky130_fd_sc_hd__xor2_1 _4735_ (.A(_3882_),
    .B(_3885_),
    .X(_3993_));
 sky130_fd_sc_hd__and2_1 _4736_ (.A(_3992_),
    .B(_3993_),
    .X(_3994_));
 sky130_fd_sc_hd__or2_1 _4737_ (.A(_3704_),
    .B(_3195_),
    .X(_3995_));
 sky130_fd_sc_hd__xnor2_1 _4738_ (.A(_3995_),
    .B(_3685_),
    .Y(_3996_));
 sky130_fd_sc_hd__xnor2_1 _4739_ (.A(_3856_),
    .B(_3880_),
    .Y(_3997_));
 sky130_fd_sc_hd__nor2_1 _4740_ (.A(_3996_),
    .B(_3997_),
    .Y(_3998_));
 sky130_fd_sc_hd__and2_1 _4741_ (.A(_3996_),
    .B(_3997_),
    .X(_3999_));
 sky130_fd_sc_hd__or2_1 _4742_ (.A(_3998_),
    .B(_3999_),
    .X(_4000_));
 sky130_fd_sc_hd__xnor2_1 _4743_ (.A(_3272_),
    .B(_3675_),
    .Y(_4001_));
 sky130_fd_sc_hd__and2_1 _4744_ (.A(_3877_),
    .B(_3878_),
    .X(_4002_));
 sky130_fd_sc_hd__or2_1 _4745_ (.A(_3879_),
    .B(_4002_),
    .X(_4003_));
 sky130_fd_sc_hd__o21ai_1 _4746_ (.A1(_3250_),
    .A2(_3327_),
    .B1(_3316_),
    .Y(_4004_));
 sky130_fd_sc_hd__xnor2_1 _4747_ (.A(_3665_),
    .B(_4004_),
    .Y(_4005_));
 sky130_fd_sc_hd__inv_2 _4748_ (.A(_4005_),
    .Y(_4006_));
 sky130_fd_sc_hd__o21a_1 _4749_ (.A1(_3876_),
    .A2(_3861_),
    .B1(_3860_),
    .X(_4007_));
 sky130_fd_sc_hd__xnor2_1 _4750_ (.A(_3875_),
    .B(_4007_),
    .Y(_4008_));
 sky130_fd_sc_hd__nor2_1 _4751_ (.A(_4006_),
    .B(_4008_),
    .Y(_4009_));
 sky130_fd_sc_hd__xnor2_1 _4752_ (.A(_3374_),
    .B(_3655_),
    .Y(_4010_));
 sky130_fd_sc_hd__xnor2_1 _4753_ (.A(_3865_),
    .B(_3874_),
    .Y(_4011_));
 sky130_fd_sc_hd__nor2_1 _4754_ (.A(_4010_),
    .B(_4011_),
    .Y(_4012_));
 sky130_fd_sc_hd__o21a_1 _4755_ (.A1(_3362_),
    .A2(_3415_),
    .B1(_3404_),
    .X(_4013_));
 sky130_fd_sc_hd__xnor2_1 _4756_ (.A(_4013_),
    .B(_3645_),
    .Y(_4014_));
 sky130_fd_sc_hd__o21a_1 _4757_ (.A1(_3863_),
    .A2(_3868_),
    .B1(_3866_),
    .X(_4015_));
 sky130_fd_sc_hd__xnor2_1 _4758_ (.A(_4015_),
    .B(_3873_),
    .Y(_4016_));
 sky130_fd_sc_hd__nor2_1 _4759_ (.A(_4014_),
    .B(_4016_),
    .Y(_4017_));
 sky130_fd_sc_hd__xnor2_1 _4760_ (.A(_3492_),
    .B(_3635_),
    .Y(_4018_));
 sky130_fd_sc_hd__a22o_1 _4761_ (.A1(_3868_),
    .A2(_3870_),
    .B1(_3869_),
    .B2(_3805_),
    .X(_4019_));
 sky130_fd_sc_hd__xnor2_1 _4762_ (.A(_3872_),
    .B(_4019_),
    .Y(_4020_));
 sky130_fd_sc_hd__nor2_1 _4763_ (.A(_4018_),
    .B(_4020_),
    .Y(_4021_));
 sky130_fd_sc_hd__a22o_1 _4764_ (.A1(_3556_),
    .A2(_3805_),
    .B1(_3809_),
    .B2(_3525_),
    .X(_4022_));
 sky130_fd_sc_hd__a22oi_1 _4765_ (.A1(_3459_),
    .A2(_2513_),
    .B1(_2425_),
    .B2(_3605_),
    .Y(_4023_));
 sky130_fd_sc_hd__or2_1 _4766_ (.A(_3626_),
    .B(_4023_),
    .X(_4024_));
 sky130_fd_sc_hd__or2_1 _4767_ (.A(_3566_),
    .B(_3616_),
    .X(_4025_));
 sky130_fd_sc_hd__xnor2_1 _4768_ (.A(_4024_),
    .B(_4025_),
    .Y(_4026_));
 sky130_fd_sc_hd__and3_1 _4769_ (.A(_3872_),
    .B(_4022_),
    .C(_4026_),
    .X(_4027_));
 sky130_fd_sc_hd__buf_2 _4770_ (.A(_3605_),
    .X(_4028_));
 sky130_fd_sc_hd__a22oi_2 _4771_ (.A1(_4028_),
    .A2(_2513_),
    .B1(_2425_),
    .B2(_3525_),
    .Y(_4029_));
 sky130_fd_sc_hd__o21ai_1 _4772_ (.A1(_3616_),
    .A2(_4029_),
    .B1(_3566_),
    .Y(_4030_));
 sky130_fd_sc_hd__o21ai_1 _4773_ (.A1(_4025_),
    .A2(_4029_),
    .B1(_4030_),
    .Y(_4031_));
 sky130_fd_sc_hd__or2b_1 _4774_ (.A(_3871_),
    .B_N(_4031_),
    .X(_4032_));
 sky130_fd_sc_hd__a21oi_1 _4775_ (.A1(_3872_),
    .A2(_4022_),
    .B1(_4026_),
    .Y(_4033_));
 sky130_fd_sc_hd__or2_1 _4776_ (.A(_4027_),
    .B(_4033_),
    .X(_4034_));
 sky130_fd_sc_hd__nor2_1 _4777_ (.A(_4032_),
    .B(_4034_),
    .Y(_4035_));
 sky130_fd_sc_hd__and2_1 _4778_ (.A(_4018_),
    .B(_4020_),
    .X(_4036_));
 sky130_fd_sc_hd__nor2_1 _4779_ (.A(_4021_),
    .B(_4036_),
    .Y(_4037_));
 sky130_fd_sc_hd__o21a_1 _4780_ (.A1(_4027_),
    .A2(_4035_),
    .B1(_4037_),
    .X(_4038_));
 sky130_fd_sc_hd__and2_1 _4781_ (.A(_4014_),
    .B(_4016_),
    .X(_4039_));
 sky130_fd_sc_hd__nor2_1 _4782_ (.A(_4017_),
    .B(_4039_),
    .Y(_4040_));
 sky130_fd_sc_hd__o21a_1 _4783_ (.A1(_4021_),
    .A2(_4038_),
    .B1(_4040_),
    .X(_4041_));
 sky130_fd_sc_hd__and2_1 _4784_ (.A(_4010_),
    .B(_4011_),
    .X(_4042_));
 sky130_fd_sc_hd__nor2_1 _4785_ (.A(_4012_),
    .B(_4042_),
    .Y(_4043_));
 sky130_fd_sc_hd__o21a_1 _4786_ (.A1(_4017_),
    .A2(_4041_),
    .B1(_4043_),
    .X(_4044_));
 sky130_fd_sc_hd__and2_1 _4787_ (.A(_4006_),
    .B(_4008_),
    .X(_4045_));
 sky130_fd_sc_hd__nor2_1 _4788_ (.A(_4009_),
    .B(_4045_),
    .Y(_4046_));
 sky130_fd_sc_hd__o21a_1 _4789_ (.A1(_4012_),
    .A2(_4044_),
    .B1(_4046_),
    .X(_4047_));
 sky130_fd_sc_hd__xor2_1 _4790_ (.A(_4001_),
    .B(_4003_),
    .X(_4048_));
 sky130_fd_sc_hd__o21ai_1 _4791_ (.A1(_4009_),
    .A2(_4047_),
    .B1(_4048_),
    .Y(_4049_));
 sky130_fd_sc_hd__o21ai_1 _4792_ (.A1(_4001_),
    .A2(_4003_),
    .B1(_4049_),
    .Y(_4050_));
 sky130_fd_sc_hd__and2b_1 _4793_ (.A_N(_4000_),
    .B(_4050_),
    .X(_4051_));
 sky130_fd_sc_hd__nor2_1 _4794_ (.A(_3992_),
    .B(_3993_),
    .Y(_4052_));
 sky130_fd_sc_hd__nor2_1 _4795_ (.A(_3994_),
    .B(_4052_),
    .Y(_4053_));
 sky130_fd_sc_hd__o21a_1 _4796_ (.A1(_3998_),
    .A2(_4051_),
    .B1(_4053_),
    .X(_4054_));
 sky130_fd_sc_hd__nand2_1 _4797_ (.A(_3988_),
    .B(_3990_),
    .Y(_4055_));
 sky130_fd_sc_hd__and2_1 _4798_ (.A(_3991_),
    .B(_4055_),
    .X(_4056_));
 sky130_fd_sc_hd__o21ai_1 _4799_ (.A1(_3994_),
    .A2(_4054_),
    .B1(_4056_),
    .Y(_4057_));
 sky130_fd_sc_hd__nor2_1 _4800_ (.A(_3984_),
    .B(_3985_),
    .Y(_4058_));
 sky130_fd_sc_hd__or2_1 _4801_ (.A(_3986_),
    .B(_4058_),
    .X(_4059_));
 sky130_fd_sc_hd__a21oi_1 _4802_ (.A1(_3991_),
    .A2(_4057_),
    .B1(_4059_),
    .Y(_4060_));
 sky130_fd_sc_hd__and2_1 _4803_ (.A(_3980_),
    .B(_3981_),
    .X(_4061_));
 sky130_fd_sc_hd__nor2_1 _4804_ (.A(_3982_),
    .B(_4061_),
    .Y(_4062_));
 sky130_fd_sc_hd__o21a_1 _4805_ (.A1(_3986_),
    .A2(_4060_),
    .B1(_4062_),
    .X(_4063_));
 sky130_fd_sc_hd__nand2_1 _4806_ (.A(_3976_),
    .B(_3977_),
    .Y(_4064_));
 sky130_fd_sc_hd__and2_1 _4807_ (.A(_3978_),
    .B(_4064_),
    .X(_4065_));
 sky130_fd_sc_hd__o21ai_1 _4808_ (.A1(_3982_),
    .A2(_4063_),
    .B1(_4065_),
    .Y(_4066_));
 sky130_fd_sc_hd__and2_1 _4809_ (.A(_3971_),
    .B(_3973_),
    .X(_4067_));
 sky130_fd_sc_hd__or2_1 _4810_ (.A(_3974_),
    .B(_4067_),
    .X(_4068_));
 sky130_fd_sc_hd__a21oi_1 _4811_ (.A1(_3978_),
    .A2(_4066_),
    .B1(_4068_),
    .Y(_4069_));
 sky130_fd_sc_hd__xnor2_1 _4812_ (.A(_3964_),
    .B(_3966_),
    .Y(_4070_));
 sky130_fd_sc_hd__o21a_1 _4813_ (.A1(_3974_),
    .A2(_4069_),
    .B1(_4070_),
    .X(_4071_));
 sky130_fd_sc_hd__or2_1 _4814_ (.A(_3959_),
    .B(_3961_),
    .X(_4072_));
 sky130_fd_sc_hd__and2_1 _4815_ (.A(_3962_),
    .B(_4072_),
    .X(_4073_));
 sky130_fd_sc_hd__o21ai_1 _4816_ (.A1(_3967_),
    .A2(_4071_),
    .B1(_4073_),
    .Y(_4074_));
 sky130_fd_sc_hd__nor2_1 _4817_ (.A(_3954_),
    .B(_3955_),
    .Y(_4075_));
 sky130_fd_sc_hd__or2_1 _4818_ (.A(_3956_),
    .B(_4075_),
    .X(_4076_));
 sky130_fd_sc_hd__a21oi_1 _4819_ (.A1(_3962_),
    .A2(_4074_),
    .B1(_4076_),
    .Y(_4077_));
 sky130_fd_sc_hd__nor2_1 _4820_ (.A(_3950_),
    .B(_3952_),
    .Y(_4078_));
 sky130_fd_sc_hd__nor2_1 _4821_ (.A(_3953_),
    .B(_4078_),
    .Y(_4079_));
 sky130_fd_sc_hd__o21a_1 _4822_ (.A1(_3956_),
    .A2(_4077_),
    .B1(_4079_),
    .X(_4080_));
 sky130_fd_sc_hd__xor2_1 _4823_ (.A(_3946_),
    .B(_3947_),
    .X(_4081_));
 sky130_fd_sc_hd__o21a_1 _4824_ (.A1(_3953_),
    .A2(_4080_),
    .B1(_4081_),
    .X(_4082_));
 sky130_fd_sc_hd__o21ba_1 _4825_ (.A1(_3946_),
    .A2(_3947_),
    .B1_N(_4082_),
    .X(_4083_));
 sky130_fd_sc_hd__o21ba_1 _4826_ (.A1(_3945_),
    .A2(_4083_),
    .B1_N(_3943_),
    .X(_4084_));
 sky130_fd_sc_hd__nor2_1 _4827_ (.A(_3937_),
    .B(_4084_),
    .Y(_4085_));
 sky130_fd_sc_hd__or2_1 _4828_ (.A(_3921_),
    .B(_3928_),
    .X(_4086_));
 sky130_fd_sc_hd__and2_1 _4829_ (.A(_3929_),
    .B(_4086_),
    .X(_4087_));
 sky130_fd_sc_hd__o21ai_1 _4830_ (.A1(_3935_),
    .A2(_4085_),
    .B1(_4087_),
    .Y(_4088_));
 sky130_fd_sc_hd__a21oi_1 _4831_ (.A1(_2458_),
    .A2(_3803_),
    .B1(_3917_),
    .Y(_4089_));
 sky130_fd_sc_hd__or2_1 _4832_ (.A(_3918_),
    .B(_4089_),
    .X(_4090_));
 sky130_fd_sc_hd__a21oi_1 _4833_ (.A1(_3929_),
    .A2(_4088_),
    .B1(_4090_),
    .Y(_4091_));
 sky130_fd_sc_hd__clkbuf_2 _4834_ (.A(_3911_),
    .X(_4092_));
 sky130_fd_sc_hd__and3_1 _4835_ (.A(_4092_),
    .B(_3808_),
    .C(_3812_),
    .X(_4093_));
 sky130_fd_sc_hd__a21oi_1 _4836_ (.A1(_4092_),
    .A2(_3808_),
    .B1(_3812_),
    .Y(_4094_));
 sky130_fd_sc_hd__or2_1 _4837_ (.A(_4093_),
    .B(_4094_),
    .X(_4095_));
 sky130_fd_sc_hd__o21ai_1 _4838_ (.A1(_3913_),
    .A2(_3915_),
    .B1(_4095_),
    .Y(_4096_));
 sky130_fd_sc_hd__o21a_1 _4839_ (.A1(_3915_),
    .A2(_4095_),
    .B1(_4096_),
    .X(_4097_));
 sky130_fd_sc_hd__nor2_1 _4840_ (.A(_3803_),
    .B(_4097_),
    .Y(_4098_));
 sky130_fd_sc_hd__and2_1 _4841_ (.A(_3803_),
    .B(_4097_),
    .X(_4099_));
 sky130_fd_sc_hd__nor2_1 _4842_ (.A(_4098_),
    .B(_4099_),
    .Y(_4100_));
 sky130_fd_sc_hd__o21a_1 _4843_ (.A1(_3918_),
    .A2(_4091_),
    .B1(_4100_),
    .X(_4101_));
 sky130_fd_sc_hd__nor3_1 _4844_ (.A(_3918_),
    .B(_4091_),
    .C(_4100_),
    .Y(_4102_));
 sky130_fd_sc_hd__nor2_1 _4845_ (.A(_4101_),
    .B(_4102_),
    .Y(_4103_));
 sky130_fd_sc_hd__buf_2 _4846_ (.A(\M1.U1.U11.u3.instance13_12.Prop_L ),
    .X(_4104_));
 sky130_fd_sc_hd__buf_2 _4847_ (.A(_4104_),
    .X(_4105_));
 sky130_fd_sc_hd__buf_2 _4848_ (.A(_4105_),
    .X(_4106_));
 sky130_fd_sc_hd__buf_2 _4849_ (.A(_4106_),
    .X(_4107_));
 sky130_fd_sc_hd__clkbuf_2 _4850_ (.A(\In2_reg[20] ),
    .X(_4108_));
 sky130_fd_sc_hd__buf_2 _4851_ (.A(_4108_),
    .X(_4109_));
 sky130_fd_sc_hd__buf_2 _4852_ (.A(_4109_),
    .X(_4110_));
 sky130_fd_sc_hd__buf_4 _4853_ (.A(_4110_),
    .X(_4111_));
 sky130_fd_sc_hd__a22o_1 _4854_ (.A1(_3819_),
    .A2(_4107_),
    .B1(_4111_),
    .B2(_3814_),
    .X(_4112_));
 sky130_fd_sc_hd__nand2_1 _4855_ (.A(_3822_),
    .B(_4106_),
    .Y(_4113_));
 sky130_fd_sc_hd__nand2_1 _4856_ (.A(_3819_),
    .B(_4111_),
    .Y(_4114_));
 sky130_fd_sc_hd__and4_1 _4857_ (.A(_3819_),
    .B(_3822_),
    .C(_4106_),
    .D(_4110_),
    .X(_4115_));
 sky130_fd_sc_hd__a21o_1 _4858_ (.A1(_4113_),
    .A2(_4114_),
    .B1(_4115_),
    .X(_4116_));
 sky130_fd_sc_hd__a22o_1 _4859_ (.A1(_3826_),
    .A2(_4106_),
    .B1(_4110_),
    .B2(_3822_),
    .X(_4117_));
 sky130_fd_sc_hd__and3_1 _4860_ (.A(_3826_),
    .B(_3828_),
    .C(_4110_),
    .X(_4118_));
 sky130_fd_sc_hd__nand2_1 _4861_ (.A(_3826_),
    .B(_4110_),
    .Y(_4119_));
 sky130_fd_sc_hd__nand2_1 _4862_ (.A(_3828_),
    .B(_4106_),
    .Y(_4120_));
 sky130_fd_sc_hd__nand2_1 _4863_ (.A(_4119_),
    .B(_4120_),
    .Y(_4121_));
 sky130_fd_sc_hd__nand2_1 _4864_ (.A(_3832_),
    .B(_4110_),
    .Y(_4122_));
 sky130_fd_sc_hd__nor2_1 _4865_ (.A(_4120_),
    .B(_4122_),
    .Y(_4123_));
 sky130_fd_sc_hd__nand2_1 _4866_ (.A(_3840_),
    .B(_4105_),
    .Y(_4124_));
 sky130_fd_sc_hd__and4_1 _4867_ (.A(_3832_),
    .B(_3840_),
    .C(_4106_),
    .D(_4110_),
    .X(_4125_));
 sky130_fd_sc_hd__a21oi_1 _4868_ (.A1(_4122_),
    .A2(_4124_),
    .B1(_4125_),
    .Y(_4126_));
 sky130_fd_sc_hd__nand2_1 _4869_ (.A(_3836_),
    .B(_4110_),
    .Y(_4127_));
 sky130_fd_sc_hd__nor2_1 _4870_ (.A(_4124_),
    .B(_4127_),
    .Y(_4128_));
 sky130_fd_sc_hd__a22o_1 _4871_ (.A1(_3844_),
    .A2(_4105_),
    .B1(_4109_),
    .B2(_3834_),
    .X(_4129_));
 sky130_fd_sc_hd__nand2_1 _4872_ (.A(_3849_),
    .B(_4105_),
    .Y(_4130_));
 sky130_fd_sc_hd__nand2_1 _4873_ (.A(_3844_),
    .B(_4109_),
    .Y(_4131_));
 sky130_fd_sc_hd__and4_1 _4874_ (.A(_3844_),
    .B(_3849_),
    .C(_4105_),
    .D(_4109_),
    .X(_4132_));
 sky130_fd_sc_hd__a21o_1 _4875_ (.A1(_4130_),
    .A2(_4131_),
    .B1(_4132_),
    .X(_4133_));
 sky130_fd_sc_hd__a22o_1 _4876_ (.A1(_3848_),
    .A2(_4105_),
    .B1(_4109_),
    .B2(_3849_),
    .X(_4134_));
 sky130_fd_sc_hd__nand2_1 _4877_ (.A(_3851_),
    .B(_4104_),
    .Y(_4135_));
 sky130_fd_sc_hd__nand2_1 _4878_ (.A(_3853_),
    .B(_4108_),
    .Y(_4136_));
 sky130_fd_sc_hd__and4_1 _4879_ (.A(_3853_),
    .B(_3857_),
    .C(_4104_),
    .D(_4108_),
    .X(_4137_));
 sky130_fd_sc_hd__a22oi_1 _4880_ (.A1(_3859_),
    .A2(_4104_),
    .B1(_4108_),
    .B2(_3857_),
    .Y(_4138_));
 sky130_fd_sc_hd__and4_1 _4881_ (.A(_3859_),
    .B(_3862_),
    .C(\M1.U1.U11.u3.instance13_12.Prop_L ),
    .D(\In2_reg[20] ),
    .X(_4139_));
 sky130_fd_sc_hd__and4_1 _4882_ (.A(_3525_),
    .B(_3556_),
    .C(\M1.U1.U11.u3.instance13_12.Prop_L ),
    .D(\In2_reg[20] ),
    .X(_4140_));
 sky130_fd_sc_hd__and2_1 _4883_ (.A(_3862_),
    .B(_4140_),
    .X(_4141_));
 sky130_fd_sc_hd__clkbuf_4 _4884_ (.A(_3525_),
    .X(_4142_));
 sky130_fd_sc_hd__and4_1 _4885_ (.A(_4028_),
    .B(_4142_),
    .C(\M1.U1.U11.u3.instance13_12.Prop_L ),
    .D(_4108_),
    .X(_4143_));
 sky130_fd_sc_hd__and4_1 _4886_ (.A(_3862_),
    .B(_4028_),
    .C(\M1.U1.U11.u3.instance13_12.Prop_L ),
    .D(\In2_reg[20] ),
    .X(_4144_));
 sky130_fd_sc_hd__a22o_1 _4887_ (.A1(_3862_),
    .A2(_4104_),
    .B1(_4108_),
    .B2(_3859_),
    .X(_4145_));
 sky130_fd_sc_hd__inv_2 _4888_ (.A(_4139_),
    .Y(_4146_));
 sky130_fd_sc_hd__o311a_1 _4889_ (.A1(_4141_),
    .A2(_4143_),
    .A3(_4144_),
    .B1(_4145_),
    .C1(_4146_),
    .X(_4147_));
 sky130_fd_sc_hd__nor2_1 _4890_ (.A(_4139_),
    .B(_4147_),
    .Y(_4148_));
 sky130_fd_sc_hd__and4_1 _4891_ (.A(_3857_),
    .B(_3859_),
    .C(_4104_),
    .D(_4108_),
    .X(_4149_));
 sky130_fd_sc_hd__o21ba_1 _4892_ (.A1(_4138_),
    .A2(_4148_),
    .B1_N(_4149_),
    .X(_4150_));
 sky130_fd_sc_hd__nand2_1 _4893_ (.A(_3857_),
    .B(_4104_),
    .Y(_4151_));
 sky130_fd_sc_hd__a21o_1 _4894_ (.A1(_4136_),
    .A2(_4151_),
    .B1(_4137_),
    .X(_4152_));
 sky130_fd_sc_hd__nor2_1 _4895_ (.A(_4150_),
    .B(_4152_),
    .Y(_4153_));
 sky130_fd_sc_hd__or2_1 _4896_ (.A(_4135_),
    .B(_4136_),
    .X(_4154_));
 sky130_fd_sc_hd__a22o_1 _4897_ (.A1(_3853_),
    .A2(_4104_),
    .B1(_4108_),
    .B2(_3851_),
    .X(_4155_));
 sky130_fd_sc_hd__o211a_1 _4898_ (.A1(_4137_),
    .A2(_4153_),
    .B1(_4154_),
    .C1(_4155_),
    .X(_4156_));
 sky130_fd_sc_hd__o21ba_1 _4899_ (.A1(_4135_),
    .A2(_4136_),
    .B1_N(_4156_),
    .X(_4157_));
 sky130_fd_sc_hd__nand2_1 _4900_ (.A(_3848_),
    .B(_4109_),
    .Y(_4158_));
 sky130_fd_sc_hd__and4_1 _4901_ (.A(_3848_),
    .B(_3851_),
    .C(_4105_),
    .D(_4109_),
    .X(_4159_));
 sky130_fd_sc_hd__a21o_1 _4902_ (.A1(_4158_),
    .A2(_4135_),
    .B1(_4159_),
    .X(_4160_));
 sky130_fd_sc_hd__o21bai_1 _4903_ (.A1(_4157_),
    .A2(_4160_),
    .B1_N(_4159_),
    .Y(_4161_));
 sky130_fd_sc_hd__o2bb2a_1 _4904_ (.A1_N(_4134_),
    .A2_N(_4161_),
    .B1(_4130_),
    .B2(_4158_),
    .X(_4162_));
 sky130_fd_sc_hd__nor2_1 _4905_ (.A(_4133_),
    .B(_4162_),
    .Y(_4163_));
 sky130_fd_sc_hd__nand2_1 _4906_ (.A(_3834_),
    .B(_4105_),
    .Y(_4164_));
 sky130_fd_sc_hd__nor2_1 _4907_ (.A(_4164_),
    .B(_4131_),
    .Y(_4165_));
 sky130_fd_sc_hd__a211o_1 _4908_ (.A1(_4129_),
    .A2(_4163_),
    .B1(_4165_),
    .C1(_4132_),
    .X(_4166_));
 sky130_fd_sc_hd__nand2_1 _4909_ (.A(_4127_),
    .B(_4164_),
    .Y(_4167_));
 sky130_fd_sc_hd__and4_1 _4910_ (.A(_3836_),
    .B(_3834_),
    .C(_4105_),
    .D(_4109_),
    .X(_4168_));
 sky130_fd_sc_hd__a21o_1 _4911_ (.A1(_4166_),
    .A2(_4167_),
    .B1(_4168_),
    .X(_4169_));
 sky130_fd_sc_hd__a22o_1 _4912_ (.A1(_3836_),
    .A2(_4106_),
    .B1(_4110_),
    .B2(_3840_),
    .X(_4170_));
 sky130_fd_sc_hd__o21a_1 _4913_ (.A1(_4128_),
    .A2(_4169_),
    .B1(_4170_),
    .X(_4171_));
 sky130_fd_sc_hd__a21o_1 _4914_ (.A1(_4126_),
    .A2(_4171_),
    .B1(_4125_),
    .X(_4172_));
 sky130_fd_sc_hd__a22oi_1 _4915_ (.A1(_3832_),
    .A2(_4106_),
    .B1(_4110_),
    .B2(_3828_),
    .Y(_4173_));
 sky130_fd_sc_hd__o21ba_1 _4916_ (.A1(_4123_),
    .A2(_4172_),
    .B1_N(_4173_),
    .X(_4174_));
 sky130_fd_sc_hd__a22o_1 _4917_ (.A1(_4106_),
    .A2(_4118_),
    .B1(_4121_),
    .B2(_4174_),
    .X(_4175_));
 sky130_fd_sc_hd__o2bb2a_1 _4918_ (.A1_N(_4117_),
    .A2_N(_4175_),
    .B1(_4113_),
    .B2(_4119_),
    .X(_4176_));
 sky130_fd_sc_hd__nor2_1 _4919_ (.A(_4116_),
    .B(_4176_),
    .Y(_4177_));
 sky130_fd_sc_hd__nand2_1 _4920_ (.A(_3814_),
    .B(_4107_),
    .Y(_4178_));
 sky130_fd_sc_hd__nor2_1 _4921_ (.A(_4178_),
    .B(_4114_),
    .Y(_4179_));
 sky130_fd_sc_hd__a211o_1 _4922_ (.A1(_4112_),
    .A2(_4177_),
    .B1(_4179_),
    .C1(_4115_),
    .X(_4180_));
 sky130_fd_sc_hd__nand2_1 _4923_ (.A(_3804_),
    .B(_4111_),
    .Y(_4181_));
 sky130_fd_sc_hd__xor2_1 _4924_ (.A(_4181_),
    .B(_4178_),
    .X(_4182_));
 sky130_fd_sc_hd__xor2_1 _4925_ (.A(_4180_),
    .B(_4182_),
    .X(_4183_));
 sky130_fd_sc_hd__buf_2 _4926_ (.A(\In2_reg[22] ),
    .X(_4184_));
 sky130_fd_sc_hd__buf_2 _4927_ (.A(_4184_),
    .X(_4185_));
 sky130_fd_sc_hd__clkbuf_2 _4928_ (.A(_4185_),
    .X(_4186_));
 sky130_fd_sc_hd__and3_1 _4929_ (.A(_3826_),
    .B(_3828_),
    .C(_4186_),
    .X(_4187_));
 sky130_fd_sc_hd__and3_1 _4930_ (.A(_3822_),
    .B(_3826_),
    .C(_4186_),
    .X(_4188_));
 sky130_fd_sc_hd__a21oi_1 _4931_ (.A1(_3822_),
    .A2(_4186_),
    .B1(_3826_),
    .Y(_4189_));
 sky130_fd_sc_hd__and3_1 _4932_ (.A(_3828_),
    .B(_3832_),
    .C(_4186_),
    .X(_4190_));
 sky130_fd_sc_hd__a21oi_1 _4933_ (.A1(_3828_),
    .A2(_4186_),
    .B1(_3832_),
    .Y(_4191_));
 sky130_fd_sc_hd__nor2_1 _4934_ (.A(_4190_),
    .B(_4191_),
    .Y(_4192_));
 sky130_fd_sc_hd__a21oi_1 _4935_ (.A1(_3832_),
    .A2(_4186_),
    .B1(_3840_),
    .Y(_4193_));
 sky130_fd_sc_hd__and3_1 _4936_ (.A(_3840_),
    .B(_3836_),
    .C(_4185_),
    .X(_4194_));
 sky130_fd_sc_hd__a21oi_1 _4937_ (.A1(_3836_),
    .A2(_4185_),
    .B1(_3834_),
    .Y(_4195_));
 sky130_fd_sc_hd__and3_1 _4938_ (.A(_3834_),
    .B(_3844_),
    .C(_4185_),
    .X(_4196_));
 sky130_fd_sc_hd__and3_1 _4939_ (.A(_3844_),
    .B(_3849_),
    .C(_4185_),
    .X(_4197_));
 sky130_fd_sc_hd__a21oi_1 _4940_ (.A1(_3844_),
    .A2(_4185_),
    .B1(_3849_),
    .Y(_4198_));
 sky130_fd_sc_hd__or2_1 _4941_ (.A(_4197_),
    .B(_4198_),
    .X(_4199_));
 sky130_fd_sc_hd__and3_1 _4942_ (.A(_3851_),
    .B(_3853_),
    .C(_4184_),
    .X(_4200_));
 sky130_fd_sc_hd__a21oi_1 _4943_ (.A1(_3851_),
    .A2(_4184_),
    .B1(_3853_),
    .Y(_4201_));
 sky130_fd_sc_hd__nor2_1 _4944_ (.A(_4200_),
    .B(_4201_),
    .Y(_4202_));
 sky130_fd_sc_hd__and3_1 _4945_ (.A(_3857_),
    .B(_3859_),
    .C(_4184_),
    .X(_4203_));
 sky130_fd_sc_hd__and3_1 _4946_ (.A(_3859_),
    .B(_3862_),
    .C(\In2_reg[22] ),
    .X(_4204_));
 sky130_fd_sc_hd__a21oi_1 _4947_ (.A1(_3859_),
    .A2(\In2_reg[22] ),
    .B1(_3862_),
    .Y(_4205_));
 sky130_fd_sc_hd__or2_1 _4948_ (.A(_4204_),
    .B(_4205_),
    .X(_4206_));
 sky130_fd_sc_hd__and3_1 _4949_ (.A(_3862_),
    .B(_4028_),
    .C(\In2_reg[22] ),
    .X(_4207_));
 sky130_fd_sc_hd__a21oi_1 _4950_ (.A1(_3862_),
    .A2(\In2_reg[22] ),
    .B1(_4028_),
    .Y(_4208_));
 sky130_fd_sc_hd__nor2_1 _4951_ (.A(_4207_),
    .B(_4208_),
    .Y(_4209_));
 sky130_fd_sc_hd__clkbuf_4 _4952_ (.A(_3556_),
    .X(_4210_));
 sky130_fd_sc_hd__o211a_1 _4953_ (.A1(_4028_),
    .A2(_4210_),
    .B1(\In2_reg[22] ),
    .C1(_4142_),
    .X(_4211_));
 sky130_fd_sc_hd__a21o_1 _4954_ (.A1(_4209_),
    .A2(_4211_),
    .B1(_4207_),
    .X(_4212_));
 sky130_fd_sc_hd__and2b_1 _4955_ (.A_N(_4206_),
    .B(_4212_),
    .X(_4213_));
 sky130_fd_sc_hd__inv_2 _4956_ (.A(_4203_),
    .Y(_4214_));
 sky130_fd_sc_hd__a21o_1 _4957_ (.A1(_3857_),
    .A2(_4184_),
    .B1(_3859_),
    .X(_4215_));
 sky130_fd_sc_hd__o211a_1 _4958_ (.A1(_4204_),
    .A2(_4213_),
    .B1(_4214_),
    .C1(_4215_),
    .X(_4216_));
 sky130_fd_sc_hd__nor2_1 _4959_ (.A(_4203_),
    .B(_4216_),
    .Y(_4217_));
 sky130_fd_sc_hd__a21oi_1 _4960_ (.A1(_3853_),
    .A2(_4184_),
    .B1(_3857_),
    .Y(_4218_));
 sky130_fd_sc_hd__and3_1 _4961_ (.A(_3853_),
    .B(_3857_),
    .C(_4184_),
    .X(_4219_));
 sky130_fd_sc_hd__o21bai_1 _4962_ (.A1(_4217_),
    .A2(_4218_),
    .B1_N(_4219_),
    .Y(_4220_));
 sky130_fd_sc_hd__a21o_1 _4963_ (.A1(_4202_),
    .A2(_4220_),
    .B1(_4200_),
    .X(_4221_));
 sky130_fd_sc_hd__a21o_1 _4964_ (.A1(_3848_),
    .A2(_4184_),
    .B1(_3851_),
    .X(_4222_));
 sky130_fd_sc_hd__a21o_1 _4965_ (.A1(_3849_),
    .A2(_4184_),
    .B1(_3848_),
    .X(_4223_));
 sky130_fd_sc_hd__nand3_1 _4966_ (.A(_3849_),
    .B(_3848_),
    .C(_4185_),
    .Y(_4224_));
 sky130_fd_sc_hd__and3_1 _4967_ (.A(_3848_),
    .B(_3851_),
    .C(_4184_),
    .X(_4225_));
 sky130_fd_sc_hd__inv_2 _4968_ (.A(_4225_),
    .Y(_4226_));
 sky130_fd_sc_hd__nand2_1 _4969_ (.A(_4224_),
    .B(_4226_),
    .Y(_4227_));
 sky130_fd_sc_hd__a31o_1 _4970_ (.A1(_4221_),
    .A2(_4222_),
    .A3(_4223_),
    .B1(_4227_),
    .X(_4228_));
 sky130_fd_sc_hd__and2b_1 _4971_ (.A_N(_4199_),
    .B(_4228_),
    .X(_4229_));
 sky130_fd_sc_hd__or2_1 _4972_ (.A(_4197_),
    .B(_4229_),
    .X(_4230_));
 sky130_fd_sc_hd__a21o_1 _4973_ (.A1(_3834_),
    .A2(_4185_),
    .B1(_3844_),
    .X(_4231_));
 sky130_fd_sc_hd__o21ai_1 _4974_ (.A1(_4196_),
    .A2(_4230_),
    .B1(_4231_),
    .Y(_4232_));
 sky130_fd_sc_hd__and3_1 _4975_ (.A(_3836_),
    .B(_3834_),
    .C(_4185_),
    .X(_4233_));
 sky130_fd_sc_hd__o21bai_1 _4976_ (.A1(_4195_),
    .A2(_4232_),
    .B1_N(_4233_),
    .Y(_4234_));
 sky130_fd_sc_hd__a21o_1 _4977_ (.A1(_3840_),
    .A2(_4185_),
    .B1(_3836_),
    .X(_4235_));
 sky130_fd_sc_hd__o21ai_1 _4978_ (.A1(_4194_),
    .A2(_4234_),
    .B1(_4235_),
    .Y(_4236_));
 sky130_fd_sc_hd__and3_1 _4979_ (.A(_3832_),
    .B(_3840_),
    .C(_4186_),
    .X(_4237_));
 sky130_fd_sc_hd__o21bai_1 _4980_ (.A1(_4193_),
    .A2(_4236_),
    .B1_N(_4237_),
    .Y(_4238_));
 sky130_fd_sc_hd__a21oi_1 _4981_ (.A1(_4192_),
    .A2(_4238_),
    .B1(_4190_),
    .Y(_4239_));
 sky130_fd_sc_hd__a21oi_1 _4982_ (.A1(_3826_),
    .A2(_4186_),
    .B1(_3828_),
    .Y(_4240_));
 sky130_fd_sc_hd__or2_1 _4983_ (.A(_4187_),
    .B(_4240_),
    .X(_4241_));
 sky130_fd_sc_hd__or3_1 _4984_ (.A(_4189_),
    .B(_4239_),
    .C(_4241_),
    .X(_4242_));
 sky130_fd_sc_hd__or3b_1 _4985_ (.A(_4187_),
    .B(_4188_),
    .C_N(_4242_),
    .X(_4243_));
 sky130_fd_sc_hd__and3_1 _4986_ (.A(_3819_),
    .B(_3822_),
    .C(_4186_),
    .X(_4244_));
 sky130_fd_sc_hd__buf_2 _4987_ (.A(_4186_),
    .X(_4245_));
 sky130_fd_sc_hd__a21o_1 _4988_ (.A1(_3819_),
    .A2(_4245_),
    .B1(_3822_),
    .X(_4246_));
 sky130_fd_sc_hd__or2b_1 _4989_ (.A(_4244_),
    .B_N(_4246_),
    .X(_4247_));
 sky130_fd_sc_hd__xnor2_1 _4990_ (.A(_4243_),
    .B(_4247_),
    .Y(_4248_));
 sky130_fd_sc_hd__xnor2_1 _4991_ (.A(_4183_),
    .B(_4248_),
    .Y(_4249_));
 sky130_fd_sc_hd__o21ai_1 _4992_ (.A1(_4178_),
    .A2(_4114_),
    .B1(_4112_),
    .Y(_4250_));
 sky130_fd_sc_hd__nor2_1 _4993_ (.A(_4115_),
    .B(_4177_),
    .Y(_4251_));
 sky130_fd_sc_hd__xnor2_1 _4994_ (.A(_4250_),
    .B(_4251_),
    .Y(_4252_));
 sky130_fd_sc_hd__nor2_1 _4995_ (.A(_4239_),
    .B(_4241_),
    .Y(_4253_));
 sky130_fd_sc_hd__nor4_1 _4996_ (.A(_4187_),
    .B(_4189_),
    .C(_4188_),
    .D(_4253_),
    .Y(_4254_));
 sky130_fd_sc_hd__o22a_1 _4997_ (.A1(_4189_),
    .A2(_4188_),
    .B1(_4253_),
    .B2(_4187_),
    .X(_4255_));
 sky130_fd_sc_hd__nor2_1 _4998_ (.A(_4254_),
    .B(_4255_),
    .Y(_4256_));
 sky130_fd_sc_hd__and2_1 _4999_ (.A(_4116_),
    .B(_4176_),
    .X(_4257_));
 sky130_fd_sc_hd__or2_1 _5000_ (.A(_4177_),
    .B(_4257_),
    .X(_4258_));
 sky130_fd_sc_hd__and2_1 _5001_ (.A(_4239_),
    .B(_4241_),
    .X(_4259_));
 sky130_fd_sc_hd__or2_1 _5002_ (.A(_4253_),
    .B(_4259_),
    .X(_4260_));
 sky130_fd_sc_hd__or2_1 _5003_ (.A(_4258_),
    .B(_4260_),
    .X(_4261_));
 sky130_fd_sc_hd__o21a_1 _5004_ (.A1(_4113_),
    .A2(_4119_),
    .B1(_4117_),
    .X(_4262_));
 sky130_fd_sc_hd__xnor2_1 _5005_ (.A(_4262_),
    .B(_4175_),
    .Y(_4263_));
 sky130_fd_sc_hd__xnor2_1 _5006_ (.A(_4192_),
    .B(_4238_),
    .Y(_4264_));
 sky130_fd_sc_hd__nor2_1 _5007_ (.A(_4263_),
    .B(_4264_),
    .Y(_4265_));
 sky130_fd_sc_hd__a22o_1 _5008_ (.A1(_4106_),
    .A2(_4118_),
    .B1(_4120_),
    .B2(_4119_),
    .X(_4266_));
 sky130_fd_sc_hd__xor2_1 _5009_ (.A(_4266_),
    .B(_4174_),
    .X(_4267_));
 sky130_fd_sc_hd__or2_1 _5010_ (.A(_4237_),
    .B(_4193_),
    .X(_4268_));
 sky130_fd_sc_hd__xnor2_1 _5011_ (.A(_4268_),
    .B(_4236_),
    .Y(_4269_));
 sky130_fd_sc_hd__nor2_1 _5012_ (.A(_4267_),
    .B(_4269_),
    .Y(_4270_));
 sky130_fd_sc_hd__and2b_1 _5013_ (.A_N(_4194_),
    .B(_4235_),
    .X(_4271_));
 sky130_fd_sc_hd__xnor2_1 _5014_ (.A(_4234_),
    .B(_4271_),
    .Y(_4272_));
 sky130_fd_sc_hd__nor2_1 _5015_ (.A(_4173_),
    .B(_4123_),
    .Y(_4273_));
 sky130_fd_sc_hd__xnor2_1 _5016_ (.A(_4172_),
    .B(_4273_),
    .Y(_4274_));
 sky130_fd_sc_hd__or2_1 _5017_ (.A(_4272_),
    .B(_4274_),
    .X(_4275_));
 sky130_fd_sc_hd__xnor2_1 _5018_ (.A(_4126_),
    .B(_4171_),
    .Y(_4276_));
 sky130_fd_sc_hd__or2_1 _5019_ (.A(_4233_),
    .B(_4195_),
    .X(_4277_));
 sky130_fd_sc_hd__xnor2_1 _5020_ (.A(_4277_),
    .B(_4232_),
    .Y(_4278_));
 sky130_fd_sc_hd__or2_1 _5021_ (.A(_4276_),
    .B(_4278_),
    .X(_4279_));
 sky130_fd_sc_hd__or2b_1 _5022_ (.A(_4196_),
    .B_N(_4231_),
    .X(_4280_));
 sky130_fd_sc_hd__xnor2_1 _5023_ (.A(_4230_),
    .B(_4280_),
    .Y(_4281_));
 sky130_fd_sc_hd__o21a_1 _5024_ (.A1(_4124_),
    .A2(_4127_),
    .B1(_4170_),
    .X(_4282_));
 sky130_fd_sc_hd__xor2_1 _5025_ (.A(_4169_),
    .B(_4282_),
    .X(_4283_));
 sky130_fd_sc_hd__nand2_1 _5026_ (.A(_4281_),
    .B(_4283_),
    .Y(_4284_));
 sky130_fd_sc_hd__or2_1 _5027_ (.A(_4281_),
    .B(_4283_),
    .X(_4285_));
 sky130_fd_sc_hd__nand2_1 _5028_ (.A(_4284_),
    .B(_4285_),
    .Y(_4286_));
 sky130_fd_sc_hd__a21o_1 _5029_ (.A1(_4127_),
    .A2(_4164_),
    .B1(_4168_),
    .X(_4287_));
 sky130_fd_sc_hd__xnor2_1 _5030_ (.A(_4166_),
    .B(_4287_),
    .Y(_4288_));
 sky130_fd_sc_hd__and2b_1 _5031_ (.A_N(_4228_),
    .B(_4199_),
    .X(_4289_));
 sky130_fd_sc_hd__nor2_1 _5032_ (.A(_4229_),
    .B(_4289_),
    .Y(_4290_));
 sky130_fd_sc_hd__o21ai_1 _5033_ (.A1(_4164_),
    .A2(_4131_),
    .B1(_4129_),
    .Y(_4291_));
 sky130_fd_sc_hd__nor2_1 _5034_ (.A(_4132_),
    .B(_4163_),
    .Y(_4292_));
 sky130_fd_sc_hd__xnor2_1 _5035_ (.A(_4291_),
    .B(_4292_),
    .Y(_4293_));
 sky130_fd_sc_hd__nand2_1 _5036_ (.A(_4223_),
    .B(_4224_),
    .Y(_4294_));
 sky130_fd_sc_hd__a21oi_1 _5037_ (.A1(_4221_),
    .A2(_4222_),
    .B1(_4225_),
    .Y(_4295_));
 sky130_fd_sc_hd__xnor2_1 _5038_ (.A(_4294_),
    .B(_4295_),
    .Y(_4296_));
 sky130_fd_sc_hd__nor2_1 _5039_ (.A(_4293_),
    .B(_4296_),
    .Y(_4297_));
 sky130_fd_sc_hd__and2_1 _5040_ (.A(_4133_),
    .B(_4162_),
    .X(_4298_));
 sky130_fd_sc_hd__or2_1 _5041_ (.A(_4163_),
    .B(_4298_),
    .X(_4299_));
 sky130_fd_sc_hd__nand2_1 _5042_ (.A(_4222_),
    .B(_4226_),
    .Y(_4300_));
 sky130_fd_sc_hd__xor2_1 _5043_ (.A(_4221_),
    .B(_4300_),
    .X(_4301_));
 sky130_fd_sc_hd__or2_1 _5044_ (.A(_4299_),
    .B(_4301_),
    .X(_4302_));
 sky130_fd_sc_hd__o21a_1 _5045_ (.A1(_4130_),
    .A2(_4158_),
    .B1(_4134_),
    .X(_4303_));
 sky130_fd_sc_hd__xnor2_1 _5046_ (.A(_4303_),
    .B(_4161_),
    .Y(_4304_));
 sky130_fd_sc_hd__xnor2_1 _5047_ (.A(_4202_),
    .B(_4220_),
    .Y(_4305_));
 sky130_fd_sc_hd__nor2_1 _5048_ (.A(_4304_),
    .B(_4305_),
    .Y(_4306_));
 sky130_fd_sc_hd__xnor2_1 _5049_ (.A(_4157_),
    .B(_4160_),
    .Y(_4307_));
 sky130_fd_sc_hd__or2_1 _5050_ (.A(_4219_),
    .B(_4218_),
    .X(_4308_));
 sky130_fd_sc_hd__xor2_1 _5051_ (.A(_4217_),
    .B(_4308_),
    .X(_4309_));
 sky130_fd_sc_hd__and2b_1 _5052_ (.A_N(_4307_),
    .B(_4309_),
    .X(_4310_));
 sky130_fd_sc_hd__a211oi_1 _5053_ (.A1(_4154_),
    .A2(_4155_),
    .B1(_4137_),
    .C1(_4153_),
    .Y(_4311_));
 sky130_fd_sc_hd__or2_1 _5054_ (.A(_4156_),
    .B(_4311_),
    .X(_4312_));
 sky130_fd_sc_hd__a211oi_1 _5055_ (.A1(_4214_),
    .A2(_4215_),
    .B1(_4204_),
    .C1(_4213_),
    .Y(_4313_));
 sky130_fd_sc_hd__or2_1 _5056_ (.A(_4216_),
    .B(_4313_),
    .X(_4314_));
 sky130_fd_sc_hd__nor2_1 _5057_ (.A(_4312_),
    .B(_4314_),
    .Y(_4315_));
 sky130_fd_sc_hd__and2_1 _5058_ (.A(_4312_),
    .B(_4314_),
    .X(_4316_));
 sky130_fd_sc_hd__nor2_1 _5059_ (.A(_4315_),
    .B(_4316_),
    .Y(_4317_));
 sky130_fd_sc_hd__xor2_1 _5060_ (.A(_4150_),
    .B(_4152_),
    .X(_4318_));
 sky130_fd_sc_hd__xnor2_1 _5061_ (.A(_4212_),
    .B(_4206_),
    .Y(_4319_));
 sky130_fd_sc_hd__xnor2_1 _5062_ (.A(_4318_),
    .B(_4319_),
    .Y(_4320_));
 sky130_fd_sc_hd__or2_1 _5063_ (.A(_4149_),
    .B(_4138_),
    .X(_4321_));
 sky130_fd_sc_hd__xnor2_1 _5064_ (.A(_4321_),
    .B(_4148_),
    .Y(_4322_));
 sky130_fd_sc_hd__xnor2_1 _5065_ (.A(_4209_),
    .B(_4211_),
    .Y(_4323_));
 sky130_fd_sc_hd__a2111oi_1 _5066_ (.A1(_4146_),
    .A2(_4145_),
    .B1(_4141_),
    .C1(_4143_),
    .D1(_4144_),
    .Y(_0096_));
 sky130_fd_sc_hd__or2_1 _5067_ (.A(_4147_),
    .B(_0096_),
    .X(_0097_));
 sky130_fd_sc_hd__nand2_2 _5068_ (.A(_3556_),
    .B(\In2_reg[22] ),
    .Y(_0098_));
 sky130_fd_sc_hd__a22o_1 _5069_ (.A1(_4028_),
    .A2(\In2_reg[22] ),
    .B1(_0098_),
    .B2(_4142_),
    .X(_0099_));
 sky130_fd_sc_hd__nand4_1 _5070_ (.A(_4028_),
    .B(_4142_),
    .C(\In2_reg[22] ),
    .D(_0098_),
    .Y(_0100_));
 sky130_fd_sc_hd__nand2_1 _5071_ (.A(_0099_),
    .B(_0100_),
    .Y(_0101_));
 sky130_fd_sc_hd__nor2_1 _5072_ (.A(_0097_),
    .B(_0101_),
    .Y(_0102_));
 sky130_fd_sc_hd__a21o_1 _5073_ (.A1(_4142_),
    .A2(\In2_reg[22] ),
    .B1(_4210_),
    .X(_0103_));
 sky130_fd_sc_hd__o21ai_1 _5074_ (.A1(_3867_),
    .A2(_0098_),
    .B1(_0103_),
    .Y(_0104_));
 sky130_fd_sc_hd__a22oi_1 _5075_ (.A1(_4028_),
    .A2(_4104_),
    .B1(_4108_),
    .B2(_3862_),
    .Y(_0105_));
 sky130_fd_sc_hd__o22a_1 _5076_ (.A1(_4140_),
    .A2(_4143_),
    .B1(_4144_),
    .B2(_0105_),
    .X(_0106_));
 sky130_fd_sc_hd__or4_1 _5077_ (.A(_4140_),
    .B(_4143_),
    .C(_4144_),
    .D(_0105_),
    .X(_0107_));
 sky130_fd_sc_hd__and2b_1 _5078_ (.A_N(_0106_),
    .B(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__or2_1 _5079_ (.A(_0104_),
    .B(_0108_),
    .X(_0109_));
 sky130_fd_sc_hd__xnor2_1 _5080_ (.A(_0104_),
    .B(_0108_),
    .Y(_0110_));
 sky130_fd_sc_hd__a22oi_1 _5081_ (.A1(_4142_),
    .A2(_4104_),
    .B1(_4108_),
    .B2(_4028_),
    .Y(_0111_));
 sky130_fd_sc_hd__nor2_1 _5082_ (.A(_4143_),
    .B(_0111_),
    .Y(_0112_));
 sky130_fd_sc_hd__xnor2_1 _5083_ (.A(_4140_),
    .B(_0112_),
    .Y(_0113_));
 sky130_fd_sc_hd__or3_1 _5084_ (.A(_0098_),
    .B(_0110_),
    .C(_0113_),
    .X(_0114_));
 sky130_fd_sc_hd__and2_1 _5085_ (.A(_0097_),
    .B(_0101_),
    .X(_0115_));
 sky130_fd_sc_hd__or2_1 _5086_ (.A(_0102_),
    .B(_0115_),
    .X(_0116_));
 sky130_fd_sc_hd__a21oi_1 _5087_ (.A1(_0109_),
    .A2(_0114_),
    .B1(_0116_),
    .Y(_0117_));
 sky130_fd_sc_hd__xor2_1 _5088_ (.A(_4322_),
    .B(_4323_),
    .X(_0118_));
 sky130_fd_sc_hd__o21a_1 _5089_ (.A1(_0102_),
    .A2(_0117_),
    .B1(_0118_),
    .X(_0119_));
 sky130_fd_sc_hd__o21ba_1 _5090_ (.A1(_4322_),
    .A2(_4323_),
    .B1_N(_0119_),
    .X(_0120_));
 sky130_fd_sc_hd__nor2_1 _5091_ (.A(_4320_),
    .B(_0120_),
    .Y(_0121_));
 sky130_fd_sc_hd__a21o_1 _5092_ (.A1(_4318_),
    .A2(_4319_),
    .B1(_0121_),
    .X(_0122_));
 sky130_fd_sc_hd__a21oi_1 _5093_ (.A1(_4317_),
    .A2(_0122_),
    .B1(_4315_),
    .Y(_0123_));
 sky130_fd_sc_hd__xnor2_1 _5094_ (.A(_4307_),
    .B(_4309_),
    .Y(_0124_));
 sky130_fd_sc_hd__and2b_1 _5095_ (.A_N(_0123_),
    .B(_0124_),
    .X(_0125_));
 sky130_fd_sc_hd__and2_1 _5096_ (.A(_4304_),
    .B(_4305_),
    .X(_0126_));
 sky130_fd_sc_hd__nor2_1 _5097_ (.A(_4306_),
    .B(_0126_),
    .Y(_0127_));
 sky130_fd_sc_hd__o21a_1 _5098_ (.A1(_4310_),
    .A2(_0125_),
    .B1(_0127_),
    .X(_0128_));
 sky130_fd_sc_hd__nand2_1 _5099_ (.A(_4299_),
    .B(_4301_),
    .Y(_0129_));
 sky130_fd_sc_hd__and2_1 _5100_ (.A(_4302_),
    .B(_0129_),
    .X(_0130_));
 sky130_fd_sc_hd__o21ai_1 _5101_ (.A1(_4306_),
    .A2(_0128_),
    .B1(_0130_),
    .Y(_0131_));
 sky130_fd_sc_hd__and2_1 _5102_ (.A(_4293_),
    .B(_4296_),
    .X(_0132_));
 sky130_fd_sc_hd__or2_1 _5103_ (.A(_4297_),
    .B(_0132_),
    .X(_0133_));
 sky130_fd_sc_hd__a21oi_1 _5104_ (.A1(_4302_),
    .A2(_0131_),
    .B1(_0133_),
    .Y(_0134_));
 sky130_fd_sc_hd__xor2_1 _5105_ (.A(_4288_),
    .B(_4290_),
    .X(_0135_));
 sky130_fd_sc_hd__o21a_1 _5106_ (.A1(_4297_),
    .A2(_0134_),
    .B1(_0135_),
    .X(_0136_));
 sky130_fd_sc_hd__a21oi_1 _5107_ (.A1(_4288_),
    .A2(_4290_),
    .B1(_0136_),
    .Y(_0137_));
 sky130_fd_sc_hd__or2_1 _5108_ (.A(_4286_),
    .B(_0137_),
    .X(_0138_));
 sky130_fd_sc_hd__nand2_1 _5109_ (.A(_4276_),
    .B(_4278_),
    .Y(_0139_));
 sky130_fd_sc_hd__nand2_1 _5110_ (.A(_4279_),
    .B(_0139_),
    .Y(_0140_));
 sky130_fd_sc_hd__a21o_1 _5111_ (.A1(_4284_),
    .A2(_0138_),
    .B1(_0140_),
    .X(_0141_));
 sky130_fd_sc_hd__nand2_1 _5112_ (.A(_4272_),
    .B(_4274_),
    .Y(_0142_));
 sky130_fd_sc_hd__nand2_1 _5113_ (.A(_4275_),
    .B(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__a21o_1 _5114_ (.A1(_4279_),
    .A2(_0141_),
    .B1(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__and2_1 _5115_ (.A(_4267_),
    .B(_4269_),
    .X(_0145_));
 sky130_fd_sc_hd__or2_1 _5116_ (.A(_4270_),
    .B(_0145_),
    .X(_0146_));
 sky130_fd_sc_hd__a21oi_1 _5117_ (.A1(_4275_),
    .A2(_0144_),
    .B1(_0146_),
    .Y(_0147_));
 sky130_fd_sc_hd__and2_1 _5118_ (.A(_4263_),
    .B(_4264_),
    .X(_0148_));
 sky130_fd_sc_hd__nor2_1 _5119_ (.A(_4265_),
    .B(_0148_),
    .Y(_0149_));
 sky130_fd_sc_hd__o21a_1 _5120_ (.A1(_4270_),
    .A2(_0147_),
    .B1(_0149_),
    .X(_0150_));
 sky130_fd_sc_hd__nand2_1 _5121_ (.A(_4258_),
    .B(_4260_),
    .Y(_0151_));
 sky130_fd_sc_hd__and2_1 _5122_ (.A(_4261_),
    .B(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__o21ai_1 _5123_ (.A1(_4265_),
    .A2(_0150_),
    .B1(_0152_),
    .Y(_0153_));
 sky130_fd_sc_hd__xnor2_1 _5124_ (.A(_4252_),
    .B(_4256_),
    .Y(_0154_));
 sky130_fd_sc_hd__a21oi_1 _5125_ (.A1(_4261_),
    .A2(_0153_),
    .B1(_0154_),
    .Y(_0155_));
 sky130_fd_sc_hd__o21bai_1 _5126_ (.A1(_4252_),
    .A2(_4256_),
    .B1_N(_0155_),
    .Y(_0156_));
 sky130_fd_sc_hd__and2b_1 _5127_ (.A_N(_4249_),
    .B(_0156_),
    .X(_0157_));
 sky130_fd_sc_hd__a21o_1 _5128_ (.A1(_4183_),
    .A2(_4248_),
    .B1(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__a2bb2o_1 _5129_ (.A1_N(_4181_),
    .A2_N(_4178_),
    .B1(_4180_),
    .B2(_4182_),
    .X(_0159_));
 sky130_fd_sc_hd__and4_1 _5130_ (.A(_3907_),
    .B(_3804_),
    .C(_4107_),
    .D(_4111_),
    .X(_0160_));
 sky130_fd_sc_hd__a22oi_1 _5131_ (.A1(_3804_),
    .A2(_4107_),
    .B1(_4111_),
    .B2(_3907_),
    .Y(_0161_));
 sky130_fd_sc_hd__or2_1 _5132_ (.A(_0160_),
    .B(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__xnor2_1 _5133_ (.A(_0159_),
    .B(_0162_),
    .Y(_0163_));
 sky130_fd_sc_hd__a21o_1 _5134_ (.A1(_4243_),
    .A2(_4246_),
    .B1(_4244_),
    .X(_0164_));
 sky130_fd_sc_hd__and3_1 _5135_ (.A(_3819_),
    .B(_3814_),
    .C(_4245_),
    .X(_0165_));
 sky130_fd_sc_hd__a21o_1 _5136_ (.A1(_3814_),
    .A2(_4245_),
    .B1(_3819_),
    .X(_0166_));
 sky130_fd_sc_hd__or2b_1 _5137_ (.A(_0165_),
    .B_N(_0166_),
    .X(_0167_));
 sky130_fd_sc_hd__xnor2_1 _5138_ (.A(_0164_),
    .B(_0167_),
    .Y(_0168_));
 sky130_fd_sc_hd__and2_1 _5139_ (.A(_0163_),
    .B(_0168_),
    .X(_0169_));
 sky130_fd_sc_hd__nor2_1 _5140_ (.A(_0163_),
    .B(_0168_),
    .Y(_0170_));
 sky130_fd_sc_hd__or2_1 _5141_ (.A(_0169_),
    .B(_0170_),
    .X(_0171_));
 sky130_fd_sc_hd__xnor2_1 _5142_ (.A(_0158_),
    .B(_0171_),
    .Y(_0172_));
 sky130_fd_sc_hd__nand2_1 _5143_ (.A(_4103_),
    .B(_0172_),
    .Y(_0173_));
 sky130_fd_sc_hd__and3_1 _5144_ (.A(_3929_),
    .B(_4088_),
    .C(_4090_),
    .X(_0174_));
 sky130_fd_sc_hd__nor2_1 _5145_ (.A(_4091_),
    .B(_0174_),
    .Y(_0175_));
 sky130_fd_sc_hd__xnor2_1 _5146_ (.A(_0156_),
    .B(_4249_),
    .Y(_0176_));
 sky130_fd_sc_hd__nand2_1 _5147_ (.A(_0175_),
    .B(_0176_),
    .Y(_0177_));
 sky130_fd_sc_hd__or2_1 _5148_ (.A(_0175_),
    .B(_0176_),
    .X(_0178_));
 sky130_fd_sc_hd__nand2_1 _5149_ (.A(_0177_),
    .B(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__or3_1 _5150_ (.A(_3935_),
    .B(_4085_),
    .C(_4087_),
    .X(_0180_));
 sky130_fd_sc_hd__and2_1 _5151_ (.A(_4088_),
    .B(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__and3_1 _5152_ (.A(_4261_),
    .B(_0153_),
    .C(_0154_),
    .X(_0182_));
 sky130_fd_sc_hd__nor2_1 _5153_ (.A(_0155_),
    .B(_0182_),
    .Y(_0183_));
 sky130_fd_sc_hd__and2_1 _5154_ (.A(_3937_),
    .B(_4084_),
    .X(_0184_));
 sky130_fd_sc_hd__or3_1 _5155_ (.A(_0152_),
    .B(_4265_),
    .C(_0150_),
    .X(_0185_));
 sky130_fd_sc_hd__and2_1 _5156_ (.A(_0153_),
    .B(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__or3b_1 _5157_ (.A(_4085_),
    .B(_0184_),
    .C_N(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__xnor2_1 _5158_ (.A(_3945_),
    .B(_4083_),
    .Y(_0188_));
 sky130_fd_sc_hd__nor3_1 _5159_ (.A(_0149_),
    .B(_4270_),
    .C(_0147_),
    .Y(_0189_));
 sky130_fd_sc_hd__or3_1 _5160_ (.A(_0150_),
    .B(_0188_),
    .C(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__nor3_1 _5161_ (.A(_4081_),
    .B(_3953_),
    .C(_4080_),
    .Y(_0191_));
 sky130_fd_sc_hd__or2_1 _5162_ (.A(_4082_),
    .B(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__and3_1 _5163_ (.A(_0146_),
    .B(_4275_),
    .C(_0144_),
    .X(_0193_));
 sky130_fd_sc_hd__or2_1 _5164_ (.A(_0147_),
    .B(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__nor2_1 _5165_ (.A(_0192_),
    .B(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__and2_1 _5166_ (.A(_0192_),
    .B(_0194_),
    .X(_0196_));
 sky130_fd_sc_hd__or2_1 _5167_ (.A(_0195_),
    .B(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__nor3_1 _5168_ (.A(_4079_),
    .B(_3956_),
    .C(_4077_),
    .Y(_0198_));
 sky130_fd_sc_hd__or2_1 _5169_ (.A(_4080_),
    .B(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__nand3_1 _5170_ (.A(_0143_),
    .B(_4279_),
    .C(_0141_),
    .Y(_0200_));
 sky130_fd_sc_hd__nand2_1 _5171_ (.A(_0144_),
    .B(_0200_),
    .Y(_0201_));
 sky130_fd_sc_hd__and3_1 _5172_ (.A(_4076_),
    .B(_3962_),
    .C(_4074_),
    .X(_0202_));
 sky130_fd_sc_hd__or2_1 _5173_ (.A(_4077_),
    .B(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__nand3_1 _5174_ (.A(_0140_),
    .B(_4284_),
    .C(_0138_),
    .Y(_0204_));
 sky130_fd_sc_hd__nand2_1 _5175_ (.A(_0141_),
    .B(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__nor2_1 _5176_ (.A(_0203_),
    .B(_0205_),
    .Y(_0206_));
 sky130_fd_sc_hd__or3_1 _5177_ (.A(_4073_),
    .B(_3967_),
    .C(_4071_),
    .X(_0207_));
 sky130_fd_sc_hd__nand2_1 _5178_ (.A(_4074_),
    .B(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__nand2_1 _5179_ (.A(_4286_),
    .B(_0137_),
    .Y(_0209_));
 sky130_fd_sc_hd__nand2_1 _5180_ (.A(_0138_),
    .B(_0209_),
    .Y(_0210_));
 sky130_fd_sc_hd__nor2_1 _5181_ (.A(_0208_),
    .B(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__nor3_1 _5182_ (.A(_4070_),
    .B(_3974_),
    .C(_4069_),
    .Y(_0212_));
 sky130_fd_sc_hd__or2_1 _5183_ (.A(_4071_),
    .B(_0212_),
    .X(_0213_));
 sky130_fd_sc_hd__nor3_1 _5184_ (.A(_0135_),
    .B(_4297_),
    .C(_0134_),
    .Y(_0214_));
 sky130_fd_sc_hd__or2_1 _5185_ (.A(_0136_),
    .B(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__nor2_1 _5186_ (.A(_0213_),
    .B(_0215_),
    .Y(_0216_));
 sky130_fd_sc_hd__and3_1 _5187_ (.A(_4068_),
    .B(_3978_),
    .C(_4066_),
    .X(_0217_));
 sky130_fd_sc_hd__or2_1 _5188_ (.A(_4069_),
    .B(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__and3_1 _5189_ (.A(_0133_),
    .B(_4302_),
    .C(_0131_),
    .X(_0219_));
 sky130_fd_sc_hd__or2_1 _5190_ (.A(_0134_),
    .B(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__nor2_1 _5191_ (.A(_0218_),
    .B(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__or3_1 _5192_ (.A(_4065_),
    .B(_3982_),
    .C(_4063_),
    .X(_0222_));
 sky130_fd_sc_hd__and2_1 _5193_ (.A(_4066_),
    .B(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__or3_1 _5194_ (.A(_0130_),
    .B(_4306_),
    .C(_0128_),
    .X(_0224_));
 sky130_fd_sc_hd__and2_1 _5195_ (.A(_0131_),
    .B(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__nand2_1 _5196_ (.A(_0223_),
    .B(_0225_),
    .Y(_0226_));
 sky130_fd_sc_hd__nor3_1 _5197_ (.A(_4062_),
    .B(_3986_),
    .C(_4060_),
    .Y(_0227_));
 sky130_fd_sc_hd__nor2_1 _5198_ (.A(_4063_),
    .B(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__nor3_1 _5199_ (.A(_0127_),
    .B(_4310_),
    .C(_0125_),
    .Y(_0229_));
 sky130_fd_sc_hd__nor2_1 _5200_ (.A(_0128_),
    .B(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__nand2_1 _5201_ (.A(_0228_),
    .B(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__and3_1 _5202_ (.A(_4059_),
    .B(_3991_),
    .C(_4057_),
    .X(_0232_));
 sky130_fd_sc_hd__or2_1 _5203_ (.A(_4060_),
    .B(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__and2b_1 _5204_ (.A_N(_0124_),
    .B(_0123_),
    .X(_0234_));
 sky130_fd_sc_hd__or2_1 _5205_ (.A(_0125_),
    .B(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__or2_1 _5206_ (.A(_0233_),
    .B(_0235_),
    .X(_0236_));
 sky130_fd_sc_hd__or3_1 _5207_ (.A(_4056_),
    .B(_3994_),
    .C(_4054_),
    .X(_0237_));
 sky130_fd_sc_hd__nand2_1 _5208_ (.A(_4057_),
    .B(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__xnor2_1 _5209_ (.A(_4317_),
    .B(_0122_),
    .Y(_0239_));
 sky130_fd_sc_hd__nor2_1 _5210_ (.A(_0238_),
    .B(_0239_),
    .Y(_0240_));
 sky130_fd_sc_hd__nor3_1 _5211_ (.A(_4053_),
    .B(_3998_),
    .C(_4051_),
    .Y(_0241_));
 sky130_fd_sc_hd__nor2_1 _5212_ (.A(_4054_),
    .B(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__and2_1 _5213_ (.A(_4320_),
    .B(_0120_),
    .X(_0243_));
 sky130_fd_sc_hd__nor2_1 _5214_ (.A(_0121_),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__and2_1 _5215_ (.A(_0242_),
    .B(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__xor2_1 _5216_ (.A(_4000_),
    .B(_4050_),
    .X(_0246_));
 sky130_fd_sc_hd__nor3_1 _5217_ (.A(_0118_),
    .B(_0102_),
    .C(_0117_),
    .Y(_0247_));
 sky130_fd_sc_hd__or3_1 _5218_ (.A(_0119_),
    .B(_0246_),
    .C(_0247_),
    .X(_0248_));
 sky130_fd_sc_hd__or3_1 _5219_ (.A(_4009_),
    .B(_4047_),
    .C(_4048_),
    .X(_0249_));
 sky130_fd_sc_hd__nand2_1 _5220_ (.A(_4049_),
    .B(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__and3_1 _5221_ (.A(_0116_),
    .B(_0109_),
    .C(_0114_),
    .X(_0251_));
 sky130_fd_sc_hd__or2_1 _5222_ (.A(_0117_),
    .B(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__nor2_1 _5223_ (.A(_0250_),
    .B(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__nor3_1 _5224_ (.A(_4012_),
    .B(_4044_),
    .C(_4046_),
    .Y(_0254_));
 sky130_fd_sc_hd__or2_1 _5225_ (.A(_4047_),
    .B(_0254_),
    .X(_0255_));
 sky130_fd_sc_hd__nor2_1 _5226_ (.A(_0098_),
    .B(_0113_),
    .Y(_0256_));
 sky130_fd_sc_hd__xnor2_1 _5227_ (.A(_0110_),
    .B(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__and2b_1 _5228_ (.A_N(_0255_),
    .B(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__nor3_1 _5229_ (.A(_4043_),
    .B(_4017_),
    .C(_4041_),
    .Y(_0259_));
 sky130_fd_sc_hd__or2_1 _5230_ (.A(_4044_),
    .B(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__and2_1 _5231_ (.A(_0098_),
    .B(_0113_),
    .X(_0261_));
 sky130_fd_sc_hd__or2_1 _5232_ (.A(_0256_),
    .B(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__nor2_1 _5233_ (.A(_0260_),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__nor3_1 _5234_ (.A(_4027_),
    .B(_4035_),
    .C(_4037_),
    .Y(_0264_));
 sky130_fd_sc_hd__nor2_1 _5235_ (.A(_4038_),
    .B(_0264_),
    .Y(_0265_));
 sky130_fd_sc_hd__and3_1 _5236_ (.A(_4210_),
    .B(_4109_),
    .C(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__nor3_1 _5237_ (.A(_4040_),
    .B(_4021_),
    .C(_4038_),
    .Y(_0267_));
 sky130_fd_sc_hd__nor2_1 _5238_ (.A(_4041_),
    .B(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__a22oi_1 _5239_ (.A1(_4210_),
    .A2(_4105_),
    .B1(_4109_),
    .B2(_4142_),
    .Y(_0269_));
 sky130_fd_sc_hd__nor2_1 _5240_ (.A(_4140_),
    .B(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__xnor2_1 _5241_ (.A(_0268_),
    .B(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__inv_2 _5242_ (.A(_0271_),
    .Y(_0272_));
 sky130_fd_sc_hd__and2_1 _5243_ (.A(_0268_),
    .B(_0270_),
    .X(_0273_));
 sky130_fd_sc_hd__a21oi_1 _5244_ (.A1(_0266_),
    .A2(_0272_),
    .B1(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__and2_1 _5245_ (.A(_0260_),
    .B(_0262_),
    .X(_0275_));
 sky130_fd_sc_hd__or2_1 _5246_ (.A(_0263_),
    .B(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__nor2_1 _5247_ (.A(_0274_),
    .B(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__xnor2_1 _5248_ (.A(_0255_),
    .B(_0257_),
    .Y(_0278_));
 sky130_fd_sc_hd__o21ai_1 _5249_ (.A1(_0263_),
    .A2(_0277_),
    .B1(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__or2b_1 _5250_ (.A(_0258_),
    .B_N(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__and2_1 _5251_ (.A(_0250_),
    .B(_0252_),
    .X(_0281_));
 sky130_fd_sc_hd__nor2_1 _5252_ (.A(_0253_),
    .B(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__and2_1 _5253_ (.A(_0280_),
    .B(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__nor2_1 _5254_ (.A(_0119_),
    .B(_0247_),
    .Y(_0284_));
 sky130_fd_sc_hd__xnor2_1 _5255_ (.A(_0246_),
    .B(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__o21ai_1 _5256_ (.A1(_0253_),
    .A2(_0283_),
    .B1(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__nor2_1 _5257_ (.A(_0242_),
    .B(_0244_),
    .Y(_0287_));
 sky130_fd_sc_hd__or2_1 _5258_ (.A(_0245_),
    .B(_0287_),
    .X(_0288_));
 sky130_fd_sc_hd__a21oi_1 _5259_ (.A1(_0248_),
    .A2(_0286_),
    .B1(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__and2_1 _5260_ (.A(_0238_),
    .B(_0239_),
    .X(_0290_));
 sky130_fd_sc_hd__nor2_1 _5261_ (.A(_0240_),
    .B(_0290_),
    .Y(_0291_));
 sky130_fd_sc_hd__o21a_1 _5262_ (.A1(_0245_),
    .A2(_0289_),
    .B1(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__nand2_1 _5263_ (.A(_0233_),
    .B(_0235_),
    .Y(_0293_));
 sky130_fd_sc_hd__and2_1 _5264_ (.A(_0236_),
    .B(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__o21ai_1 _5265_ (.A1(_0240_),
    .A2(_0292_),
    .B1(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__or2_1 _5266_ (.A(_0228_),
    .B(_0230_),
    .X(_0296_));
 sky130_fd_sc_hd__nand2_1 _5267_ (.A(_0231_),
    .B(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__a21o_1 _5268_ (.A1(_0236_),
    .A2(_0295_),
    .B1(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__or2_1 _5269_ (.A(_0223_),
    .B(_0225_),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_1 _5270_ (.A(_0226_),
    .B(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__a21o_1 _5271_ (.A1(_0231_),
    .A2(_0298_),
    .B1(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__and2_1 _5272_ (.A(_0218_),
    .B(_0220_),
    .X(_0302_));
 sky130_fd_sc_hd__or2_1 _5273_ (.A(_0221_),
    .B(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__a21oi_1 _5274_ (.A1(_0226_),
    .A2(_0301_),
    .B1(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__and2_1 _5275_ (.A(_0213_),
    .B(_0215_),
    .X(_0305_));
 sky130_fd_sc_hd__or2_1 _5276_ (.A(_0216_),
    .B(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__o21ba_1 _5277_ (.A1(_0221_),
    .A2(_0304_),
    .B1_N(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__and2_1 _5278_ (.A(_0208_),
    .B(_0210_),
    .X(_0308_));
 sky130_fd_sc_hd__nor2_1 _5279_ (.A(_0211_),
    .B(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__o21a_1 _5280_ (.A1(_0216_),
    .A2(_0307_),
    .B1(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__and2_1 _5281_ (.A(_0203_),
    .B(_0205_),
    .X(_0311_));
 sky130_fd_sc_hd__nor2_1 _5282_ (.A(_0206_),
    .B(_0311_),
    .Y(_0312_));
 sky130_fd_sc_hd__o21a_1 _5283_ (.A1(_0211_),
    .A2(_0310_),
    .B1(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__xor2_1 _5284_ (.A(_0199_),
    .B(_0201_),
    .X(_0314_));
 sky130_fd_sc_hd__o21a_1 _5285_ (.A1(_0206_),
    .A2(_0313_),
    .B1(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__o21bai_2 _5286_ (.A1(_0199_),
    .A2(_0201_),
    .B1_N(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__and2b_1 _5287_ (.A_N(_0197_),
    .B(_0316_),
    .X(_0317_));
 sky130_fd_sc_hd__nor2_1 _5288_ (.A(_0150_),
    .B(_0189_),
    .Y(_0318_));
 sky130_fd_sc_hd__xnor2_1 _5289_ (.A(_0188_),
    .B(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__o21ai_1 _5290_ (.A1(_0195_),
    .A2(_0317_),
    .B1(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__or2_1 _5291_ (.A(_4085_),
    .B(_0184_),
    .X(_0321_));
 sky130_fd_sc_hd__xor2_1 _5292_ (.A(_0321_),
    .B(_0186_),
    .X(_0322_));
 sky130_fd_sc_hd__a21o_1 _5293_ (.A1(_0190_),
    .A2(_0320_),
    .B1(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__xnor2_1 _5294_ (.A(_0181_),
    .B(_0183_),
    .Y(_0324_));
 sky130_fd_sc_hd__a21o_1 _5295_ (.A1(_0187_),
    .A2(_0323_),
    .B1(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__a21bo_1 _5296_ (.A1(_0181_),
    .A2(_0183_),
    .B1_N(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__nand2b_1 _5297_ (.A_N(_0179_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__or2_1 _5298_ (.A(_4103_),
    .B(_0172_),
    .X(_0328_));
 sky130_fd_sc_hd__nand2_1 _5299_ (.A(_0173_),
    .B(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__a21o_1 _5300_ (.A1(_0177_),
    .A2(_0327_),
    .B1(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__nand2_1 _5301_ (.A(_0173_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__nor2_1 _5302_ (.A(_3915_),
    .B(_4093_),
    .Y(_0332_));
 sky130_fd_sc_hd__and2_1 _5303_ (.A(_3808_),
    .B(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__o21ai_1 _5304_ (.A1(_4098_),
    .A2(_4101_),
    .B1(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__or3_1 _5305_ (.A(_4098_),
    .B(_4101_),
    .C(_0333_),
    .X(_0335_));
 sky130_fd_sc_hd__and2_1 _5306_ (.A(_0334_),
    .B(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__and2b_1 _5307_ (.A_N(_0171_),
    .B(_0158_),
    .X(_0337_));
 sky130_fd_sc_hd__and2b_1 _5308_ (.A_N(_0162_),
    .B(_0159_),
    .X(_0338_));
 sky130_fd_sc_hd__nand4_1 _5309_ (.A(_4092_),
    .B(_3907_),
    .C(_4107_),
    .D(_4111_),
    .Y(_0339_));
 sky130_fd_sc_hd__a22o_1 _5310_ (.A1(_3907_),
    .A2(_4107_),
    .B1(_4111_),
    .B2(_4092_),
    .X(_0340_));
 sky130_fd_sc_hd__o211a_1 _5311_ (.A1(_0160_),
    .A2(_0338_),
    .B1(_0339_),
    .C1(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__a211o_1 _5312_ (.A1(_0339_),
    .A2(_0340_),
    .B1(_0160_),
    .C1(_0338_),
    .X(_0342_));
 sky130_fd_sc_hd__and2b_1 _5313_ (.A_N(_0341_),
    .B(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__a21oi_1 _5314_ (.A1(_0164_),
    .A2(_0166_),
    .B1(_0165_),
    .Y(_0344_));
 sky130_fd_sc_hd__and3_1 _5315_ (.A(_3804_),
    .B(_3814_),
    .C(_4245_),
    .X(_0345_));
 sky130_fd_sc_hd__a21oi_1 _5316_ (.A1(_3804_),
    .A2(_4245_),
    .B1(_3814_),
    .Y(_0346_));
 sky130_fd_sc_hd__or2_1 _5317_ (.A(_0345_),
    .B(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__xor2_1 _5318_ (.A(_0344_),
    .B(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__and2_1 _5319_ (.A(_0343_),
    .B(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__nor2_1 _5320_ (.A(_0343_),
    .B(_0348_),
    .Y(_0350_));
 sky130_fd_sc_hd__nor2_1 _5321_ (.A(_0349_),
    .B(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__o21a_1 _5322_ (.A1(_0169_),
    .A2(_0337_),
    .B1(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__nor3_1 _5323_ (.A(_0169_),
    .B(_0337_),
    .C(_0351_),
    .Y(_0353_));
 sky130_fd_sc_hd__nor2_1 _5324_ (.A(_0352_),
    .B(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__nand2_1 _5325_ (.A(_0336_),
    .B(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__or2_1 _5326_ (.A(_0336_),
    .B(_0354_),
    .X(_0356_));
 sky130_fd_sc_hd__nand2_1 _5327_ (.A(_0355_),
    .B(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__xnor2_2 _5328_ (.A(_0331_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__buf_2 _5329_ (.A(\M1.U1.U8.u3.instance7_6.Prop_L ),
    .X(_0359_));
 sky130_fd_sc_hd__buf_2 _5330_ (.A(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__buf_2 _5331_ (.A(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_2 _5332_ (.A(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__buf_2 _5333_ (.A(\In2_reg[14] ),
    .X(_0363_));
 sky130_fd_sc_hd__buf_2 _5334_ (.A(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__buf_2 _5335_ (.A(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__buf_2 _5336_ (.A(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__and4_1 _5337_ (.A(_2579_),
    .B(_2634_),
    .C(_0362_),
    .D(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__nand2_1 _5338_ (.A(_2579_),
    .B(_0362_),
    .Y(_0368_));
 sky130_fd_sc_hd__nand2_1 _5339_ (.A(_2491_),
    .B(_0366_),
    .Y(_0369_));
 sky130_fd_sc_hd__nor2_1 _5340_ (.A(_0368_),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__and2_1 _5341_ (.A(_0368_),
    .B(_0369_),
    .X(_0371_));
 sky130_fd_sc_hd__a22o_1 _5342_ (.A1(_2733_),
    .A2(_0361_),
    .B1(_0366_),
    .B2(_2689_),
    .X(_0372_));
 sky130_fd_sc_hd__and4_1 _5343_ (.A(_2722_),
    .B(_2788_),
    .C(_0361_),
    .D(_0365_),
    .X(_0373_));
 sky130_fd_sc_hd__and4_1 _5344_ (.A(_2799_),
    .B(_2843_),
    .C(_0361_),
    .D(_0365_),
    .X(_0374_));
 sky130_fd_sc_hd__a22oi_1 _5345_ (.A1(_2799_),
    .A2(_0361_),
    .B1(_0365_),
    .B2(_2733_),
    .Y(_0375_));
 sky130_fd_sc_hd__or2_1 _5346_ (.A(_0373_),
    .B(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__a22oi_1 _5347_ (.A1(_2843_),
    .A2(_0361_),
    .B1(_0365_),
    .B2(_2799_),
    .Y(_0377_));
 sky130_fd_sc_hd__or2_1 _5348_ (.A(_0374_),
    .B(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__and4_1 _5349_ (.A(_2843_),
    .B(_2876_),
    .C(_0361_),
    .D(_0365_),
    .X(_0379_));
 sky130_fd_sc_hd__a22oi_1 _5350_ (.A1(_2876_),
    .A2(_0361_),
    .B1(_0365_),
    .B2(_2843_),
    .Y(_0380_));
 sky130_fd_sc_hd__nor2_1 _5351_ (.A(_0379_),
    .B(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__a22o_1 _5352_ (.A1(_2997_),
    .A2(_0360_),
    .B1(_0365_),
    .B2(_2920_),
    .X(_0382_));
 sky130_fd_sc_hd__and4_1 _5353_ (.A(_2997_),
    .B(_3041_),
    .C(_0360_),
    .D(_0364_),
    .X(_0383_));
 sky130_fd_sc_hd__nand2_1 _5354_ (.A(_3041_),
    .B(_0360_),
    .Y(_0384_));
 sky130_fd_sc_hd__nand2_1 _5355_ (.A(_3096_),
    .B(_0364_),
    .Y(_0385_));
 sky130_fd_sc_hd__nor2_1 _5356_ (.A(_0384_),
    .B(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__and4_1 _5357_ (.A(_3096_),
    .B(_3140_),
    .C(_0360_),
    .D(_0364_),
    .X(_0387_));
 sky130_fd_sc_hd__nand2_1 _5358_ (.A(_3140_),
    .B(_0360_),
    .Y(_0388_));
 sky130_fd_sc_hd__a21oi_1 _5359_ (.A1(_0385_),
    .A2(_0388_),
    .B1(_0387_),
    .Y(_0389_));
 sky130_fd_sc_hd__a22o_1 _5360_ (.A1(_3184_),
    .A2(_0360_),
    .B1(_0364_),
    .B2(_3140_),
    .X(_0390_));
 sky130_fd_sc_hd__nand2_1 _5361_ (.A(_3239_),
    .B(_0360_),
    .Y(_0391_));
 sky130_fd_sc_hd__nand2_1 _5362_ (.A(_3184_),
    .B(_0364_),
    .Y(_0392_));
 sky130_fd_sc_hd__and4_1 _5363_ (.A(_3184_),
    .B(_3239_),
    .C(_0359_),
    .D(_0364_),
    .X(_0393_));
 sky130_fd_sc_hd__a21o_1 _5364_ (.A1(_0391_),
    .A2(_0392_),
    .B1(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__a22o_1 _5365_ (.A1(_3305_),
    .A2(_0359_),
    .B1(_0363_),
    .B2(_3239_),
    .X(_0395_));
 sky130_fd_sc_hd__and3_1 _5366_ (.A(_3305_),
    .B(_3355_),
    .C(_0359_),
    .X(_0396_));
 sky130_fd_sc_hd__nand2_1 _5367_ (.A(_3305_),
    .B(_0363_),
    .Y(_0397_));
 sky130_fd_sc_hd__nand2_1 _5368_ (.A(_3355_),
    .B(_0359_),
    .Y(_0398_));
 sky130_fd_sc_hd__a22o_1 _5369_ (.A1(_0397_),
    .A2(_0398_),
    .B1(_0396_),
    .B2(_0363_),
    .X(_0399_));
 sky130_fd_sc_hd__nand2_1 _5370_ (.A(_3393_),
    .B(_0363_),
    .Y(_0400_));
 sky130_fd_sc_hd__nor2_1 _5371_ (.A(_0398_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__nand2_1 _5372_ (.A(_3459_),
    .B(_0359_),
    .Y(_0402_));
 sky130_fd_sc_hd__and4_1 _5373_ (.A(_3387_),
    .B(_3459_),
    .C(_0359_),
    .D(_0363_),
    .X(_0403_));
 sky130_fd_sc_hd__a21oi_1 _5374_ (.A1(_0400_),
    .A2(_0402_),
    .B1(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__and4_1 _5375_ (.A(_3596_),
    .B(_3514_),
    .C(\M1.U1.U8.u3.instance7_6.Prop_L ),
    .D(\In2_reg[14] ),
    .X(_0405_));
 sky130_fd_sc_hd__a22oi_1 _5376_ (.A1(_3605_),
    .A2(_0359_),
    .B1(_0363_),
    .B2(_3448_),
    .Y(_0406_));
 sky130_fd_sc_hd__nand2_1 _5377_ (.A(_3596_),
    .B(_0363_),
    .Y(_0407_));
 sky130_fd_sc_hd__nand2_1 _5378_ (.A(_3514_),
    .B(\M1.U1.U8.u3.instance7_6.Prop_L ),
    .Y(_0408_));
 sky130_fd_sc_hd__a21o_1 _5379_ (.A1(_0407_),
    .A2(_0408_),
    .B1(_0405_),
    .X(_0409_));
 sky130_fd_sc_hd__nand2_1 _5380_ (.A(_3546_),
    .B(\In2_reg[14] ),
    .Y(_0410_));
 sky130_fd_sc_hd__or2_2 _5381_ (.A(_0408_),
    .B(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__nor3_1 _5382_ (.A(_0406_),
    .B(_0409_),
    .C(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__nor2_1 _5383_ (.A(_0402_),
    .B(_0407_),
    .Y(_0413_));
 sky130_fd_sc_hd__or3_1 _5384_ (.A(_0405_),
    .B(_0412_),
    .C(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__a21o_1 _5385_ (.A1(_0404_),
    .A2(_0414_),
    .B1(_0403_),
    .X(_0415_));
 sky130_fd_sc_hd__a22o_1 _5386_ (.A1(_3393_),
    .A2(_0359_),
    .B1(_0363_),
    .B2(_3355_),
    .X(_0416_));
 sky130_fd_sc_hd__o21a_1 _5387_ (.A1(_0401_),
    .A2(_0415_),
    .B1(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__nor2b_1 _5388_ (.A(_0399_),
    .B_N(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__a21o_1 _5389_ (.A1(_0364_),
    .A2(_0396_),
    .B1(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__o2bb2a_1 _5390_ (.A1_N(_0395_),
    .A2_N(_0419_),
    .B1(_0391_),
    .B2(_0397_),
    .X(_0420_));
 sky130_fd_sc_hd__nor2_1 _5391_ (.A(_0394_),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__nor2_1 _5392_ (.A(_0388_),
    .B(_0392_),
    .Y(_0422_));
 sky130_fd_sc_hd__a211o_1 _5393_ (.A1(_0390_),
    .A2(_0421_),
    .B1(_0422_),
    .C1(_0393_),
    .X(_0423_));
 sky130_fd_sc_hd__and2_1 _5394_ (.A(_0389_),
    .B(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__or2_1 _5395_ (.A(_0384_),
    .B(_0385_),
    .X(_0425_));
 sky130_fd_sc_hd__a22o_1 _5396_ (.A1(_3096_),
    .A2(_0360_),
    .B1(_0364_),
    .B2(_3041_),
    .X(_0426_));
 sky130_fd_sc_hd__o211a_1 _5397_ (.A1(_0387_),
    .A2(_0424_),
    .B1(_0425_),
    .C1(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_1 _5398_ (.A(_2997_),
    .B(_0364_),
    .Y(_0428_));
 sky130_fd_sc_hd__a21oi_1 _5399_ (.A1(_0428_),
    .A2(_0384_),
    .B1(_0383_),
    .Y(_0429_));
 sky130_fd_sc_hd__o21a_1 _5400_ (.A1(_0386_),
    .A2(_0427_),
    .B1(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__or2_1 _5401_ (.A(_0383_),
    .B(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__nand2_1 _5402_ (.A(_2920_),
    .B(_0360_),
    .Y(_0432_));
 sky130_fd_sc_hd__o2bb2a_1 _5403_ (.A1_N(_0382_),
    .A2_N(_0431_),
    .B1(_0432_),
    .B2(_0428_),
    .X(_0433_));
 sky130_fd_sc_hd__nand2_1 _5404_ (.A(_2876_),
    .B(_0365_),
    .Y(_0434_));
 sky130_fd_sc_hd__and4_1 _5405_ (.A(_2876_),
    .B(_2920_),
    .C(_0361_),
    .D(_0365_),
    .X(_0435_));
 sky130_fd_sc_hd__a21o_1 _5406_ (.A1(_0432_),
    .A2(_0434_),
    .B1(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__o21bai_2 _5407_ (.A1(_0433_),
    .A2(_0436_),
    .B1_N(_0435_),
    .Y(_0437_));
 sky130_fd_sc_hd__a21oi_2 _5408_ (.A1(_0437_),
    .A2(_0381_),
    .B1(_0379_),
    .Y(_0438_));
 sky130_fd_sc_hd__nor3_1 _5409_ (.A(_0376_),
    .B(_0378_),
    .C(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__or3_1 _5410_ (.A(_0373_),
    .B(_0374_),
    .C(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__nand4_1 _5411_ (.A(_2689_),
    .B(_2733_),
    .C(_0361_),
    .D(_0366_),
    .Y(_0441_));
 sky130_fd_sc_hd__a21bo_1 _5412_ (.A1(_0372_),
    .A2(_0440_),
    .B1_N(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__and4_1 _5413_ (.A(_2689_),
    .B(_2634_),
    .C(_0362_),
    .D(_0366_),
    .X(_0443_));
 sky130_fd_sc_hd__a22o_1 _5414_ (.A1(_2689_),
    .A2(_0362_),
    .B1(_0366_),
    .B2(_2634_),
    .X(_0444_));
 sky130_fd_sc_hd__o21a_1 _5415_ (.A1(_0442_),
    .A2(_0443_),
    .B1(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__a22oi_1 _5416_ (.A1(_3814_),
    .A2(_0362_),
    .B1(_0366_),
    .B2(_2579_),
    .Y(_0446_));
 sky130_fd_sc_hd__nor2_1 _5417_ (.A(_0367_),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__and2_1 _5418_ (.A(_0445_),
    .B(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__and2b_1 _5419_ (.A_N(_0371_),
    .B(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__or3_1 _5420_ (.A(_0367_),
    .B(_0370_),
    .C(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__nand2_1 _5421_ (.A(_3911_),
    .B(_0362_),
    .Y(_0451_));
 sky130_fd_sc_hd__a22o_1 _5422_ (.A1(_2491_),
    .A2(_0362_),
    .B1(_0366_),
    .B2(_3911_),
    .X(_0452_));
 sky130_fd_sc_hd__o21a_1 _5423_ (.A1(_0369_),
    .A2(_0451_),
    .B1(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__and2_1 _5424_ (.A(_0450_),
    .B(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__and3_1 _5425_ (.A(_3911_),
    .B(_0362_),
    .C(_0366_),
    .X(_0455_));
 sky130_fd_sc_hd__nor2_1 _5426_ (.A(_0454_),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__buf_2 _5427_ (.A(\In2_reg[12] ),
    .X(_0457_));
 sky130_fd_sc_hd__buf_2 _5428_ (.A(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__buf_2 _5429_ (.A(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__buf_2 _5430_ (.A(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__nand2_1 _5431_ (.A(_0460_),
    .B(_2579_),
    .Y(_0461_));
 sky130_fd_sc_hd__buf_2 _5432_ (.A(\M1.U1.U7.u3.instance5_4.Prop_L ),
    .X(_0462_));
 sky130_fd_sc_hd__buf_2 _5433_ (.A(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__buf_2 _5434_ (.A(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__buf_2 _5435_ (.A(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__nand2_1 _5436_ (.A(_2634_),
    .B(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__and4_1 _5437_ (.A(_0460_),
    .B(_2568_),
    .C(_2634_),
    .D(_0465_),
    .X(_0467_));
 sky130_fd_sc_hd__a21o_1 _5438_ (.A1(_0461_),
    .A2(_0466_),
    .B1(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__nand2_1 _5439_ (.A(_2689_),
    .B(_0460_),
    .Y(_0469_));
 sky130_fd_sc_hd__a22o_1 _5440_ (.A1(_0460_),
    .A2(_2623_),
    .B1(_0464_),
    .B2(_2678_),
    .X(_0470_));
 sky130_fd_sc_hd__o21ai_1 _5441_ (.A1(_0466_),
    .A2(_0469_),
    .B1(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__nand2_1 _5442_ (.A(_2722_),
    .B(_0464_),
    .Y(_0472_));
 sky130_fd_sc_hd__and4_1 _5443_ (.A(_2678_),
    .B(_2733_),
    .C(_0459_),
    .D(_0464_),
    .X(_0473_));
 sky130_fd_sc_hd__a21o_1 _5444_ (.A1(_0469_),
    .A2(_0472_),
    .B1(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__or2_1 _5445_ (.A(_0471_),
    .B(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__nand2_1 _5446_ (.A(_2788_),
    .B(_0459_),
    .Y(_0476_));
 sky130_fd_sc_hd__a22o_1 _5447_ (.A1(_2722_),
    .A2(_0459_),
    .B1(_0464_),
    .B2(_2799_),
    .X(_0477_));
 sky130_fd_sc_hd__o21a_1 _5448_ (.A1(_0472_),
    .A2(_0476_),
    .B1(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__a22o_1 _5449_ (.A1(_2832_),
    .A2(_0459_),
    .B1(_0464_),
    .B2(_2865_),
    .X(_0479_));
 sky130_fd_sc_hd__and4_1 _5450_ (.A(_2865_),
    .B(_2920_),
    .C(_0459_),
    .D(_0464_),
    .X(_0480_));
 sky130_fd_sc_hd__nand2_1 _5451_ (.A(_2909_),
    .B(_0463_),
    .Y(_0481_));
 sky130_fd_sc_hd__nand2_1 _5452_ (.A(_2986_),
    .B(_0459_),
    .Y(_0482_));
 sky130_fd_sc_hd__nor2_1 _5453_ (.A(_0481_),
    .B(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__and4_1 _5454_ (.A(_2986_),
    .B(_3041_),
    .C(_0458_),
    .D(_0463_),
    .X(_0484_));
 sky130_fd_sc_hd__nand2_1 _5455_ (.A(_3030_),
    .B(_0463_),
    .Y(_0485_));
 sky130_fd_sc_hd__a21oi_1 _5456_ (.A1(_0482_),
    .A2(_0485_),
    .B1(_0484_),
    .Y(_0486_));
 sky130_fd_sc_hd__a22o_1 _5457_ (.A1(_3030_),
    .A2(_0458_),
    .B1(_0463_),
    .B2(_3096_),
    .X(_0487_));
 sky130_fd_sc_hd__nand2_1 _5458_ (.A(_3140_),
    .B(_0463_),
    .Y(_0488_));
 sky130_fd_sc_hd__nand2_1 _5459_ (.A(_3085_),
    .B(_0458_),
    .Y(_0489_));
 sky130_fd_sc_hd__and4_1 _5460_ (.A(_3085_),
    .B(_3129_),
    .C(_0458_),
    .D(_0463_),
    .X(_0490_));
 sky130_fd_sc_hd__a21o_1 _5461_ (.A1(_0488_),
    .A2(_0489_),
    .B1(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__a22o_1 _5462_ (.A1(_3129_),
    .A2(_0458_),
    .B1(_0463_),
    .B2(_3184_),
    .X(_0492_));
 sky130_fd_sc_hd__nand2_1 _5463_ (.A(_3173_),
    .B(_0458_),
    .Y(_0493_));
 sky130_fd_sc_hd__nand2_1 _5464_ (.A(_3239_),
    .B(_0463_),
    .Y(_0494_));
 sky130_fd_sc_hd__and4_1 _5465_ (.A(_3173_),
    .B(_3239_),
    .C(_0458_),
    .D(_0462_),
    .X(_0495_));
 sky130_fd_sc_hd__a21oi_1 _5466_ (.A1(_0493_),
    .A2(_0494_),
    .B1(_0495_),
    .Y(_0496_));
 sky130_fd_sc_hd__and2_1 _5467_ (.A(_3305_),
    .B(_0462_),
    .X(_0497_));
 sky130_fd_sc_hd__a21o_1 _5468_ (.A1(_3239_),
    .A2(_0457_),
    .B1(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__and4_1 _5469_ (.A(_3228_),
    .B(_3305_),
    .C(_0457_),
    .D(_0462_),
    .X(_0499_));
 sky130_fd_sc_hd__and2_1 _5470_ (.A(_3349_),
    .B(_0457_),
    .X(_0500_));
 sky130_fd_sc_hd__a22o_1 _5471_ (.A1(_3294_),
    .A2(_0457_),
    .B1(_0462_),
    .B2(_3355_),
    .X(_0501_));
 sky130_fd_sc_hd__and3_1 _5472_ (.A(_3387_),
    .B(_0462_),
    .C(_0500_),
    .X(_0502_));
 sky130_fd_sc_hd__a22o_1 _5473_ (.A1(_3387_),
    .A2(_0457_),
    .B1(_0462_),
    .B2(_3448_),
    .X(_0503_));
 sky130_fd_sc_hd__and4_2 _5474_ (.A(_3514_),
    .B(_3546_),
    .C(\In2_reg[12] ),
    .D(\M1.U1.U7.u3.instance5_4.Prop_L ),
    .X(_0504_));
 sky130_fd_sc_hd__and4_1 _5475_ (.A(_3596_),
    .B(_3503_),
    .C(\In2_reg[12] ),
    .D(\M1.U1.U7.u3.instance5_4.Prop_L ),
    .X(_0505_));
 sky130_fd_sc_hd__and4_1 _5476_ (.A(_3448_),
    .B(_3596_),
    .C(_0457_),
    .D(\M1.U1.U7.u3.instance5_4.Prop_L ),
    .X(_0506_));
 sky130_fd_sc_hd__a211o_1 _5477_ (.A1(_3448_),
    .A2(_0504_),
    .B1(_0505_),
    .C1(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__and4_1 _5478_ (.A(_3387_),
    .B(_3448_),
    .C(_0457_),
    .D(\M1.U1.U7.u3.instance5_4.Prop_L ),
    .X(_0508_));
 sky130_fd_sc_hd__a21o_1 _5479_ (.A1(_0503_),
    .A2(_0507_),
    .B1(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__a21o_1 _5480_ (.A1(_3393_),
    .A2(_0462_),
    .B1(_0500_),
    .X(_0510_));
 sky130_fd_sc_hd__o21a_1 _5481_ (.A1(_0502_),
    .A2(_0509_),
    .B1(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__a22o_1 _5482_ (.A1(_0497_),
    .A2(_0500_),
    .B1(_0501_),
    .B2(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__or2_1 _5483_ (.A(_0499_),
    .B(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__a31o_1 _5484_ (.A1(_0496_),
    .A2(_0498_),
    .A3(_0513_),
    .B1(_0495_),
    .X(_0514_));
 sky130_fd_sc_hd__o2bb2a_1 _5485_ (.A1_N(_0492_),
    .A2_N(_0514_),
    .B1(_0488_),
    .B2(_0493_),
    .X(_0515_));
 sky130_fd_sc_hd__nor2_1 _5486_ (.A(_0491_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__nor2_1 _5487_ (.A(_0485_),
    .B(_0489_),
    .Y(_0517_));
 sky130_fd_sc_hd__a211o_1 _5488_ (.A1(_0487_),
    .A2(_0516_),
    .B1(_0517_),
    .C1(_0490_),
    .X(_0518_));
 sky130_fd_sc_hd__and2_1 _5489_ (.A(_0486_),
    .B(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__or2_1 _5490_ (.A(_0481_),
    .B(_0482_),
    .X(_0520_));
 sky130_fd_sc_hd__a22o_1 _5491_ (.A1(_2920_),
    .A2(_0459_),
    .B1(_0464_),
    .B2(_2997_),
    .X(_0521_));
 sky130_fd_sc_hd__o211a_1 _5492_ (.A1(_0484_),
    .A2(_0519_),
    .B1(_0520_),
    .C1(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__nand2_1 _5493_ (.A(_2865_),
    .B(_0459_),
    .Y(_0523_));
 sky130_fd_sc_hd__a21oi_1 _5494_ (.A1(_0523_),
    .A2(_0481_),
    .B1(_0480_),
    .Y(_0524_));
 sky130_fd_sc_hd__o21a_1 _5495_ (.A1(_0483_),
    .A2(_0522_),
    .B1(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__or2_1 _5496_ (.A(_0480_),
    .B(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__nand2_1 _5497_ (.A(_2832_),
    .B(_0464_),
    .Y(_0527_));
 sky130_fd_sc_hd__o2bb2a_1 _5498_ (.A1_N(_0479_),
    .A2_N(_0526_),
    .B1(_0527_),
    .B2(_0523_),
    .X(_0528_));
 sky130_fd_sc_hd__and4_1 _5499_ (.A(_2788_),
    .B(_2832_),
    .C(_0459_),
    .D(_0464_),
    .X(_0529_));
 sky130_fd_sc_hd__a21o_1 _5500_ (.A1(_0527_),
    .A2(_0476_),
    .B1(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__o21bai_2 _5501_ (.A1(_0528_),
    .A2(_0530_),
    .B1_N(_0529_),
    .Y(_0531_));
 sky130_fd_sc_hd__nor2_1 _5502_ (.A(_0472_),
    .B(_0476_),
    .Y(_0532_));
 sky130_fd_sc_hd__a21oi_2 _5503_ (.A1(_0478_),
    .A2(_0531_),
    .B1(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__o21bai_1 _5504_ (.A1(_0466_),
    .A2(_0469_),
    .B1_N(_0473_),
    .Y(_0534_));
 sky130_fd_sc_hd__o21ba_1 _5505_ (.A1(_0475_),
    .A2(_0533_),
    .B1_N(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__o21bai_2 _5506_ (.A1(_0468_),
    .A2(_0535_),
    .B1_N(_0467_),
    .Y(_0536_));
 sky130_fd_sc_hd__and4_1 _5507_ (.A(_0460_),
    .B(_2480_),
    .C(_2579_),
    .D(_0465_),
    .X(_0537_));
 sky130_fd_sc_hd__a22o_1 _5508_ (.A1(_0460_),
    .A2(_2480_),
    .B1(_2579_),
    .B2(_0465_),
    .X(_0538_));
 sky130_fd_sc_hd__o21ai_2 _5509_ (.A1(_0536_),
    .A2(_0537_),
    .B1(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__a22o_1 _5510_ (.A1(_0460_),
    .A2(_3801_),
    .B1(_2491_),
    .B2(_0465_),
    .X(_0540_));
 sky130_fd_sc_hd__nand4_1 _5511_ (.A(_0460_),
    .B(_3801_),
    .C(_2491_),
    .D(_0465_),
    .Y(_0541_));
 sky130_fd_sc_hd__nand2_1 _5512_ (.A(_0540_),
    .B(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__nor2_1 _5513_ (.A(_0539_),
    .B(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__and3_1 _5514_ (.A(_0460_),
    .B(_3801_),
    .C(_0465_),
    .X(_0544_));
 sky130_fd_sc_hd__nor2_1 _5515_ (.A(_0543_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__a21oi_1 _5516_ (.A1(_3911_),
    .A2(_0362_),
    .B1(_0366_),
    .Y(_0546_));
 sky130_fd_sc_hd__o21a_1 _5517_ (.A1(_0455_),
    .A2(_0546_),
    .B1(_0369_),
    .X(_0547_));
 sky130_fd_sc_hd__nor2_1 _5518_ (.A(_0455_),
    .B(_0546_),
    .Y(_0548_));
 sky130_fd_sc_hd__mux2_1 _5519_ (.A0(_0547_),
    .A1(_0548_),
    .S(_0454_),
    .X(_0549_));
 sky130_fd_sc_hd__nor2_1 _5520_ (.A(_0545_),
    .B(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__xor2_1 _5521_ (.A(_0450_),
    .B(_0453_),
    .X(_0551_));
 sky130_fd_sc_hd__and3_1 _5522_ (.A(_0465_),
    .B(_0545_),
    .C(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__a21oi_1 _5523_ (.A1(_0465_),
    .A2(_0545_),
    .B1(_0551_),
    .Y(_0553_));
 sky130_fd_sc_hd__or2_1 _5524_ (.A(_0552_),
    .B(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__or4_1 _5525_ (.A(_0367_),
    .B(_0448_),
    .C(_0370_),
    .D(_0371_),
    .X(_0555_));
 sky130_fd_sc_hd__o22ai_1 _5526_ (.A1(_0367_),
    .A2(_0448_),
    .B1(_0370_),
    .B2(_0371_),
    .Y(_0556_));
 sky130_fd_sc_hd__nand2_1 _5527_ (.A(_0555_),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__a21oi_1 _5528_ (.A1(_3911_),
    .A2(_0465_),
    .B1(_0460_),
    .Y(_0558_));
 sky130_fd_sc_hd__or2_1 _5529_ (.A(_0544_),
    .B(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__nand2_1 _5530_ (.A(_0541_),
    .B(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__mux2_1 _5531_ (.A0(_0560_),
    .A1(_0559_),
    .S(_0543_),
    .X(_0561_));
 sky130_fd_sc_hd__and2_1 _5532_ (.A(_0557_),
    .B(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__nor2_1 _5533_ (.A(_0557_),
    .B(_0561_),
    .Y(_0563_));
 sky130_fd_sc_hd__nor2_1 _5534_ (.A(_0562_),
    .B(_0563_),
    .Y(_0564_));
 sky130_fd_sc_hd__xnor2_1 _5535_ (.A(_0539_),
    .B(_0542_),
    .Y(_0565_));
 sky130_fd_sc_hd__xnor2_1 _5536_ (.A(_0445_),
    .B(_0447_),
    .Y(_0566_));
 sky130_fd_sc_hd__and2_1 _5537_ (.A(_0536_),
    .B(_0537_),
    .X(_0567_));
 sky130_fd_sc_hd__o22a_1 _5538_ (.A1(_0538_),
    .A2(_0536_),
    .B1(_0539_),
    .B2(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__nand2_1 _5539_ (.A(_0442_),
    .B(_0443_),
    .Y(_0569_));
 sky130_fd_sc_hd__o2bb2a_1 _5540_ (.A1_N(_0445_),
    .A2_N(_0569_),
    .B1(_0444_),
    .B2(_0442_),
    .X(_0570_));
 sky130_fd_sc_hd__and2_1 _5541_ (.A(_0568_),
    .B(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__xnor2_1 _5542_ (.A(_0468_),
    .B(_0535_),
    .Y(_0572_));
 sky130_fd_sc_hd__nand2_1 _5543_ (.A(_0441_),
    .B(_0372_),
    .Y(_0573_));
 sky130_fd_sc_hd__xor2_1 _5544_ (.A(_0573_),
    .B(_0440_),
    .X(_0574_));
 sky130_fd_sc_hd__or2_1 _5545_ (.A(_0572_),
    .B(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__nand2_1 _5546_ (.A(_0572_),
    .B(_0574_),
    .Y(_0576_));
 sky130_fd_sc_hd__and2_1 _5547_ (.A(_0575_),
    .B(_0576_),
    .X(_0577_));
 sky130_fd_sc_hd__o21ba_1 _5548_ (.A1(_0474_),
    .A2(_0533_),
    .B1_N(_0473_),
    .X(_0578_));
 sky130_fd_sc_hd__xnor2_1 _5549_ (.A(_0471_),
    .B(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__o21ba_1 _5550_ (.A1(_0378_),
    .A2(_0438_),
    .B1_N(_0374_),
    .X(_0580_));
 sky130_fd_sc_hd__xnor2_1 _5551_ (.A(_0376_),
    .B(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__nand2_1 _5552_ (.A(_0579_),
    .B(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__or2_1 _5553_ (.A(_0579_),
    .B(_0581_),
    .X(_0583_));
 sky130_fd_sc_hd__xnor2_1 _5554_ (.A(_0474_),
    .B(_0533_),
    .Y(_0584_));
 sky130_fd_sc_hd__xnor2_1 _5555_ (.A(_0378_),
    .B(_0438_),
    .Y(_0585_));
 sky130_fd_sc_hd__xnor2_1 _5556_ (.A(_0478_),
    .B(_0531_),
    .Y(_0586_));
 sky130_fd_sc_hd__xnor2_1 _5557_ (.A(_0381_),
    .B(_0437_),
    .Y(_0587_));
 sky130_fd_sc_hd__xnor2_1 _5558_ (.A(_0528_),
    .B(_0530_),
    .Y(_0588_));
 sky130_fd_sc_hd__xnor2_1 _5559_ (.A(_0433_),
    .B(_0436_),
    .Y(_0589_));
 sky130_fd_sc_hd__nor2_1 _5560_ (.A(_0588_),
    .B(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__o21a_1 _5561_ (.A1(_0527_),
    .A2(_0523_),
    .B1(_0479_),
    .X(_0591_));
 sky130_fd_sc_hd__xnor2_1 _5562_ (.A(_0591_),
    .B(_0526_),
    .Y(_0592_));
 sky130_fd_sc_hd__o21a_1 _5563_ (.A1(_0432_),
    .A2(_0428_),
    .B1(_0382_),
    .X(_0593_));
 sky130_fd_sc_hd__xnor2_1 _5564_ (.A(_0593_),
    .B(_0431_),
    .Y(_0594_));
 sky130_fd_sc_hd__or2_1 _5565_ (.A(_0592_),
    .B(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__nor3_1 _5566_ (.A(_0483_),
    .B(_0522_),
    .C(_0524_),
    .Y(_0596_));
 sky130_fd_sc_hd__nor2_1 _5567_ (.A(_0525_),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__nor3_1 _5568_ (.A(_0386_),
    .B(_0427_),
    .C(_0429_),
    .Y(_0598_));
 sky130_fd_sc_hd__nor2_1 _5569_ (.A(_0430_),
    .B(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__and2_1 _5570_ (.A(_0597_),
    .B(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__a211oi_1 _5571_ (.A1(_0520_),
    .A2(_0521_),
    .B1(_0484_),
    .C1(_0519_),
    .Y(_0601_));
 sky130_fd_sc_hd__or2_1 _5572_ (.A(_0522_),
    .B(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__a211oi_1 _5573_ (.A1(_0425_),
    .A2(_0426_),
    .B1(_0387_),
    .C1(_0424_),
    .Y(_0603_));
 sky130_fd_sc_hd__or2_1 _5574_ (.A(_0427_),
    .B(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__nor2_1 _5575_ (.A(_0602_),
    .B(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__xnor2_1 _5576_ (.A(_0486_),
    .B(_0518_),
    .Y(_0606_));
 sky130_fd_sc_hd__xnor2_1 _5577_ (.A(_0389_),
    .B(_0423_),
    .Y(_0607_));
 sky130_fd_sc_hd__nor2_1 _5578_ (.A(_0606_),
    .B(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__and2_1 _5579_ (.A(_0606_),
    .B(_0607_),
    .X(_0609_));
 sky130_fd_sc_hd__or2_1 _5580_ (.A(_0608_),
    .B(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__o21ai_1 _5581_ (.A1(_0485_),
    .A2(_0489_),
    .B1(_0487_),
    .Y(_0611_));
 sky130_fd_sc_hd__nor2_1 _5582_ (.A(_0490_),
    .B(_0516_),
    .Y(_0612_));
 sky130_fd_sc_hd__xnor2_1 _5583_ (.A(_0611_),
    .B(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__o21ai_1 _5584_ (.A1(_0388_),
    .A2(_0392_),
    .B1(_0390_),
    .Y(_0614_));
 sky130_fd_sc_hd__nor2_1 _5585_ (.A(_0393_),
    .B(_0421_),
    .Y(_0615_));
 sky130_fd_sc_hd__xnor2_1 _5586_ (.A(_0614_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__xnor2_1 _5587_ (.A(_0491_),
    .B(_0515_),
    .Y(_0617_));
 sky130_fd_sc_hd__xnor2_1 _5588_ (.A(_0394_),
    .B(_0420_),
    .Y(_0618_));
 sky130_fd_sc_hd__nor2_1 _5589_ (.A(_0617_),
    .B(_0618_),
    .Y(_0619_));
 sky130_fd_sc_hd__o21a_1 _5590_ (.A1(_0488_),
    .A2(_0493_),
    .B1(_0492_),
    .X(_0620_));
 sky130_fd_sc_hd__xnor2_1 _5591_ (.A(_0620_),
    .B(_0514_),
    .Y(_0621_));
 sky130_fd_sc_hd__o21a_1 _5592_ (.A1(_0391_),
    .A2(_0397_),
    .B1(_0395_),
    .X(_0622_));
 sky130_fd_sc_hd__xnor2_1 _5593_ (.A(_0622_),
    .B(_0419_),
    .Y(_0623_));
 sky130_fd_sc_hd__nor2_1 _5594_ (.A(_0621_),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand2_1 _5595_ (.A(_0498_),
    .B(_0513_),
    .Y(_0625_));
 sky130_fd_sc_hd__xor2_1 _5596_ (.A(_0496_),
    .B(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__xor2_1 _5597_ (.A(_0399_),
    .B(_0417_),
    .X(_0627_));
 sky130_fd_sc_hd__nor2_1 _5598_ (.A(_0626_),
    .B(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__o21ai_1 _5599_ (.A1(_0398_),
    .A2(_0400_),
    .B1(_0416_),
    .Y(_0629_));
 sky130_fd_sc_hd__xnor2_1 _5600_ (.A(_0415_),
    .B(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__or2b_1 _5601_ (.A(_0499_),
    .B_N(_0498_),
    .X(_0631_));
 sky130_fd_sc_hd__xnor2_1 _5602_ (.A(_0512_),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__and2_1 _5603_ (.A(_0630_),
    .B(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__a21bo_1 _5604_ (.A1(_0497_),
    .A2(_0500_),
    .B1_N(_0501_),
    .X(_0634_));
 sky130_fd_sc_hd__xor2_1 _5605_ (.A(_0634_),
    .B(_0511_),
    .X(_0635_));
 sky130_fd_sc_hd__xnor2_1 _5606_ (.A(_0404_),
    .B(_0414_),
    .Y(_0636_));
 sky130_fd_sc_hd__nor2_1 _5607_ (.A(_0635_),
    .B(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__nor2_1 _5608_ (.A(_0406_),
    .B(_0413_),
    .Y(_0638_));
 sky130_fd_sc_hd__or2b_1 _5609_ (.A(_0405_),
    .B_N(_0411_),
    .X(_0639_));
 sky130_fd_sc_hd__xnor2_1 _5610_ (.A(_0638_),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__nor2_1 _5611_ (.A(_0510_),
    .B(_0509_),
    .Y(_0641_));
 sky130_fd_sc_hd__o2bb2a_1 _5612_ (.A1_N(_0502_),
    .A2_N(_0509_),
    .B1(_0511_),
    .B2(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__nor2_1 _5613_ (.A(_0640_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__or2b_1 _5614_ (.A(_0508_),
    .B_N(_0503_),
    .X(_0644_));
 sky130_fd_sc_hd__xor2_1 _5615_ (.A(_0644_),
    .B(_0507_),
    .X(_0645_));
 sky130_fd_sc_hd__xnor2_1 _5616_ (.A(_0409_),
    .B(_0411_),
    .Y(_0646_));
 sky130_fd_sc_hd__or2_1 _5617_ (.A(_0645_),
    .B(_0646_),
    .X(_0647_));
 sky130_fd_sc_hd__a22o_1 _5618_ (.A1(_3556_),
    .A2(_0359_),
    .B1(_0363_),
    .B2(_3525_),
    .X(_0648_));
 sky130_fd_sc_hd__a22oi_1 _5619_ (.A1(_3448_),
    .A2(_0457_),
    .B1(_0462_),
    .B2(_3605_),
    .Y(_0649_));
 sky130_fd_sc_hd__o22ai_1 _5620_ (.A1(_0504_),
    .A2(_0505_),
    .B1(_0506_),
    .B2(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__or4_1 _5621_ (.A(_0504_),
    .B(_0505_),
    .C(_0506_),
    .D(_0649_),
    .X(_0651_));
 sky130_fd_sc_hd__nand2_1 _5622_ (.A(_0650_),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__a22oi_1 _5623_ (.A1(_3605_),
    .A2(_0457_),
    .B1(_0462_),
    .B2(_3514_),
    .Y(_0653_));
 sky130_fd_sc_hd__nor2_1 _5624_ (.A(_0505_),
    .B(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__xnor2_1 _5625_ (.A(_0504_),
    .B(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__or2_1 _5626_ (.A(_0410_),
    .B(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__nand2_1 _5627_ (.A(_0411_),
    .B(_0648_),
    .Y(_0657_));
 sky130_fd_sc_hd__xor2_1 _5628_ (.A(_0657_),
    .B(_0652_),
    .X(_0658_));
 sky130_fd_sc_hd__nor2_1 _5629_ (.A(_0656_),
    .B(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__a31o_1 _5630_ (.A1(_0411_),
    .A2(_0648_),
    .A3(_0652_),
    .B1(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__nand2_1 _5631_ (.A(_0645_),
    .B(_0646_),
    .Y(_0661_));
 sky130_fd_sc_hd__and2_1 _5632_ (.A(_0647_),
    .B(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__nand2_1 _5633_ (.A(_0660_),
    .B(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__and2_1 _5634_ (.A(_0640_),
    .B(_0642_),
    .X(_0664_));
 sky130_fd_sc_hd__or2_1 _5635_ (.A(_0643_),
    .B(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__a21oi_1 _5636_ (.A1(_0647_),
    .A2(_0663_),
    .B1(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__and2_1 _5637_ (.A(_0635_),
    .B(_0636_),
    .X(_0667_));
 sky130_fd_sc_hd__nor2_1 _5638_ (.A(_0637_),
    .B(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__o21a_1 _5639_ (.A1(_0643_),
    .A2(_0666_),
    .B1(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__nor2_1 _5640_ (.A(_0630_),
    .B(_0632_),
    .Y(_0670_));
 sky130_fd_sc_hd__nor2_1 _5641_ (.A(_0633_),
    .B(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__o21a_1 _5642_ (.A1(_0637_),
    .A2(_0669_),
    .B1(_0671_),
    .X(_0672_));
 sky130_fd_sc_hd__and2_1 _5643_ (.A(_0626_),
    .B(_0627_),
    .X(_0673_));
 sky130_fd_sc_hd__nor2_1 _5644_ (.A(_0628_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__o21a_1 _5645_ (.A1(_0633_),
    .A2(_0672_),
    .B1(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__and2_1 _5646_ (.A(_0621_),
    .B(_0623_),
    .X(_0676_));
 sky130_fd_sc_hd__nor2_1 _5647_ (.A(_0624_),
    .B(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__o21a_1 _5648_ (.A1(_0628_),
    .A2(_0675_),
    .B1(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__and2_1 _5649_ (.A(_0617_),
    .B(_0618_),
    .X(_0679_));
 sky130_fd_sc_hd__nor2_1 _5650_ (.A(_0619_),
    .B(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__o21a_1 _5651_ (.A1(_0624_),
    .A2(_0678_),
    .B1(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__xor2_1 _5652_ (.A(_0613_),
    .B(_0616_),
    .X(_0682_));
 sky130_fd_sc_hd__o21a_1 _5653_ (.A1(_0619_),
    .A2(_0681_),
    .B1(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__o21bai_1 _5654_ (.A1(_0613_),
    .A2(_0616_),
    .B1_N(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__and2b_1 _5655_ (.A_N(_0610_),
    .B(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__and2_1 _5656_ (.A(_0602_),
    .B(_0604_),
    .X(_0686_));
 sky130_fd_sc_hd__nor2_1 _5657_ (.A(_0605_),
    .B(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__o21a_1 _5658_ (.A1(_0608_),
    .A2(_0685_),
    .B1(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__nor2_1 _5659_ (.A(_0597_),
    .B(_0599_),
    .Y(_0689_));
 sky130_fd_sc_hd__nor2_1 _5660_ (.A(_0600_),
    .B(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__o21a_1 _5661_ (.A1(_0605_),
    .A2(_0688_),
    .B1(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__nand2_1 _5662_ (.A(_0592_),
    .B(_0594_),
    .Y(_0692_));
 sky130_fd_sc_hd__and2_1 _5663_ (.A(_0595_),
    .B(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__o21ai_1 _5664_ (.A1(_0600_),
    .A2(_0691_),
    .B1(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__nand2_1 _5665_ (.A(_0588_),
    .B(_0589_),
    .Y(_0695_));
 sky130_fd_sc_hd__or2b_1 _5666_ (.A(_0590_),
    .B_N(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__a21oi_1 _5667_ (.A1(_0595_),
    .A2(_0694_),
    .B1(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__xor2_1 _5668_ (.A(_0586_),
    .B(_0587_),
    .X(_0698_));
 sky130_fd_sc_hd__o21ai_1 _5669_ (.A1(_0590_),
    .A2(_0697_),
    .B1(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__o21a_1 _5670_ (.A1(_0586_),
    .A2(_0587_),
    .B1(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__o21a_1 _5671_ (.A1(_0584_),
    .A2(_0585_),
    .B1(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__a21o_1 _5672_ (.A1(_0584_),
    .A2(_0585_),
    .B1(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__nand2_1 _5673_ (.A(_0583_),
    .B(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__and2_1 _5674_ (.A(_0582_),
    .B(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__nand2_1 _5675_ (.A(_0577_),
    .B(_0704_),
    .Y(_0705_));
 sky130_fd_sc_hd__nor2_1 _5676_ (.A(_0568_),
    .B(_0570_),
    .Y(_0706_));
 sky130_fd_sc_hd__or2_1 _5677_ (.A(_0571_),
    .B(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__a21oi_1 _5678_ (.A1(_0575_),
    .A2(_0705_),
    .B1(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__xor2_1 _5679_ (.A(_0565_),
    .B(_0566_),
    .X(_0709_));
 sky130_fd_sc_hd__o21ai_1 _5680_ (.A1(_0571_),
    .A2(_0708_),
    .B1(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__o21ai_1 _5681_ (.A1(_0565_),
    .A2(_0566_),
    .B1(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__a21o_1 _5682_ (.A1(_0564_),
    .A2(_0711_),
    .B1(_0562_),
    .X(_0712_));
 sky130_fd_sc_hd__and2b_1 _5683_ (.A_N(_0554_),
    .B(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__and2_1 _5684_ (.A(_0545_),
    .B(_0549_),
    .X(_0714_));
 sky130_fd_sc_hd__nor2_1 _5685_ (.A(_0550_),
    .B(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__o21a_1 _5686_ (.A1(_0552_),
    .A2(_0713_),
    .B1(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__and2_1 _5687_ (.A(_0362_),
    .B(_0456_),
    .X(_0717_));
 sky130_fd_sc_hd__o21ai_1 _5688_ (.A1(_0550_),
    .A2(_0716_),
    .B1(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__buf_2 _5689_ (.A(\M1.U1.U6.u3.instance3_2.Prop_L ),
    .X(_0719_));
 sky130_fd_sc_hd__buf_2 _5690_ (.A(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__buf_2 _5691_ (.A(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__buf_2 _5692_ (.A(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__inv_2 _5693_ (.A(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__buf_2 _5694_ (.A(\In2_reg[8] ),
    .X(_0724_));
 sky130_fd_sc_hd__buf_2 _5695_ (.A(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__buf_2 _5696_ (.A(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__clkbuf_2 _5697_ (.A(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__buf_2 _5698_ (.A(\M1.U1.U5.u3.instance1_0.Prop_L ),
    .X(_0728_));
 sky130_fd_sc_hd__buf_2 _5699_ (.A(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__buf_2 _5700_ (.A(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__clkbuf_2 _5701_ (.A(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__and4_1 _5702_ (.A(_0727_),
    .B(_0731_),
    .C(_2469_),
    .D(_2568_),
    .X(_0732_));
 sky130_fd_sc_hd__and4_1 _5703_ (.A(_0727_),
    .B(_0731_),
    .C(_2557_),
    .D(_2623_),
    .X(_0733_));
 sky130_fd_sc_hd__and4_1 _5704_ (.A(_0727_),
    .B(_2667_),
    .C(_0731_),
    .D(_2612_),
    .X(_0734_));
 sky130_fd_sc_hd__a22oi_1 _5705_ (.A1(_2667_),
    .A2(_0731_),
    .B1(_2612_),
    .B2(_0727_),
    .Y(_0735_));
 sky130_fd_sc_hd__nor2_1 _5706_ (.A(_0734_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__nand2_1 _5707_ (.A(_0727_),
    .B(_2667_),
    .Y(_0737_));
 sky130_fd_sc_hd__nand2_1 _5708_ (.A(_0730_),
    .B(_2711_),
    .Y(_0738_));
 sky130_fd_sc_hd__and4_1 _5709_ (.A(_0726_),
    .B(_0730_),
    .C(_2711_),
    .D(_2777_),
    .X(_0739_));
 sky130_fd_sc_hd__and4_1 _5710_ (.A(_0726_),
    .B(_0730_),
    .C(_2777_),
    .D(_2821_),
    .X(_0740_));
 sky130_fd_sc_hd__a22oi_1 _5711_ (.A1(_0726_),
    .A2(_2777_),
    .B1(_2821_),
    .B2(_0730_),
    .Y(_0741_));
 sky130_fd_sc_hd__nor2_1 _5712_ (.A(_0740_),
    .B(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__and4_1 _5713_ (.A(_0725_),
    .B(_0729_),
    .C(\In1_reg[14] ),
    .D(_2898_),
    .X(_0743_));
 sky130_fd_sc_hd__a22oi_1 _5714_ (.A1(_0725_),
    .A2(\In1_reg[14] ),
    .B1(_2898_),
    .B2(_0729_),
    .Y(_0744_));
 sky130_fd_sc_hd__or2_1 _5715_ (.A(_0743_),
    .B(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__and4_1 _5716_ (.A(_0725_),
    .B(_0729_),
    .C(\In1_reg[15] ),
    .D(\In1_reg[14] ),
    .X(_0746_));
 sky130_fd_sc_hd__a22oi_1 _5717_ (.A1(_0725_),
    .A2(\In1_reg[15] ),
    .B1(_2854_),
    .B2(_0729_),
    .Y(_0747_));
 sky130_fd_sc_hd__or2_1 _5718_ (.A(_0746_),
    .B(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__nor2_1 _5719_ (.A(_0745_),
    .B(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__and4_1 _5720_ (.A(_0726_),
    .B(_0729_),
    .C(_2898_),
    .D(_2975_),
    .X(_0750_));
 sky130_fd_sc_hd__a22oi_1 _5721_ (.A1(_0726_),
    .A2(_2898_),
    .B1(_2986_),
    .B2(_0730_),
    .Y(_0751_));
 sky130_fd_sc_hd__nor2_1 _5722_ (.A(_0750_),
    .B(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__nand2_1 _5723_ (.A(_0730_),
    .B(_3019_),
    .Y(_0753_));
 sky130_fd_sc_hd__nand2_1 _5724_ (.A(_0725_),
    .B(_3085_),
    .Y(_0754_));
 sky130_fd_sc_hd__a22o_1 _5725_ (.A1(_0725_),
    .A2(_3019_),
    .B1(_3085_),
    .B2(_0729_),
    .X(_0755_));
 sky130_fd_sc_hd__o21a_1 _5726_ (.A1(_0753_),
    .A2(_0754_),
    .B1(_0755_),
    .X(_0756_));
 sky130_fd_sc_hd__nand2_1 _5727_ (.A(_0729_),
    .B(_3129_),
    .Y(_0757_));
 sky130_fd_sc_hd__and4_1 _5728_ (.A(_0725_),
    .B(_0729_),
    .C(_3074_),
    .D(_3129_),
    .X(_0758_));
 sky130_fd_sc_hd__a21o_1 _5729_ (.A1(_0754_),
    .A2(_0757_),
    .B1(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__a22o_1 _5730_ (.A1(_0724_),
    .A2(_3228_),
    .B1(_3305_),
    .B2(_0728_),
    .X(_0760_));
 sky130_fd_sc_hd__nand2_1 _5731_ (.A(_0724_),
    .B(_3294_),
    .Y(_0761_));
 sky130_fd_sc_hd__nand2_1 _5732_ (.A(_0728_),
    .B(_3355_),
    .Y(_0762_));
 sky130_fd_sc_hd__and4_1 _5733_ (.A(_0724_),
    .B(_0728_),
    .C(_3294_),
    .D(_3349_),
    .X(_0763_));
 sky130_fd_sc_hd__a21o_1 _5734_ (.A1(_0761_),
    .A2(_0762_),
    .B1(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__and3_1 _5735_ (.A(_0724_),
    .B(_0728_),
    .C(_3349_),
    .X(_0765_));
 sky130_fd_sc_hd__a22o_1 _5736_ (.A1(_0724_),
    .A2(_3349_),
    .B1(_3387_),
    .B2(_0728_),
    .X(_0766_));
 sky130_fd_sc_hd__a22o_1 _5737_ (.A1(_0724_),
    .A2(_3387_),
    .B1(_3448_),
    .B2(_0728_),
    .X(_0767_));
 sky130_fd_sc_hd__a22o_1 _5738_ (.A1(\In2_reg[8] ),
    .A2(_3448_),
    .B1(_3596_),
    .B2(\M1.U1.U5.u3.instance1_0.Prop_L ),
    .X(_0768_));
 sky130_fd_sc_hd__o2111a_1 _5739_ (.A1(_3596_),
    .A2(_3546_),
    .B1(_3514_),
    .C1(\In2_reg[8] ),
    .D1(\M1.U1.U5.u3.instance1_0.Prop_L ),
    .X(_0769_));
 sky130_fd_sc_hd__and4_1 _5740_ (.A(\In2_reg[8] ),
    .B(\M1.U1.U5.u3.instance1_0.Prop_L ),
    .C(_3437_),
    .D(_3596_),
    .X(_0770_));
 sky130_fd_sc_hd__a21o_1 _5741_ (.A1(_0768_),
    .A2(_0769_),
    .B1(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__and4_1 _5742_ (.A(\In2_reg[8] ),
    .B(\M1.U1.U5.u3.instance1_0.Prop_L ),
    .C(_3387_),
    .D(_3448_),
    .X(_0772_));
 sky130_fd_sc_hd__a21o_1 _5743_ (.A1(_0767_),
    .A2(_0771_),
    .B1(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__a22oi_2 _5744_ (.A1(_3393_),
    .A2(_0765_),
    .B1(_0766_),
    .B2(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__o21bai_1 _5745_ (.A1(_0764_),
    .A2(_0774_),
    .B1_N(_0763_),
    .Y(_0775_));
 sky130_fd_sc_hd__nand2_1 _5746_ (.A(_0728_),
    .B(_3228_),
    .Y(_0776_));
 sky130_fd_sc_hd__o2bb2a_1 _5747_ (.A1_N(_0760_),
    .A2_N(_0775_),
    .B1(_0776_),
    .B2(_0761_),
    .X(_0777_));
 sky130_fd_sc_hd__nand2_1 _5748_ (.A(_0725_),
    .B(_3173_),
    .Y(_0778_));
 sky130_fd_sc_hd__and4_1 _5749_ (.A(_0724_),
    .B(_0728_),
    .C(_3173_),
    .D(_3228_),
    .X(_0779_));
 sky130_fd_sc_hd__a21oi_1 _5750_ (.A1(_0778_),
    .A2(_0776_),
    .B1(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__nor2b_1 _5751_ (.A(_0777_),
    .B_N(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__a22o_1 _5752_ (.A1(_0725_),
    .A2(_3129_),
    .B1(_3173_),
    .B2(_0729_),
    .X(_0782_));
 sky130_fd_sc_hd__o21a_1 _5753_ (.A1(_0757_),
    .A2(_0778_),
    .B1(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__o21bai_1 _5754_ (.A1(_0757_),
    .A2(_0778_),
    .B1_N(_0779_),
    .Y(_0784_));
 sky130_fd_sc_hd__a21oi_1 _5755_ (.A1(_0781_),
    .A2(_0783_),
    .B1(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__nor2_1 _5756_ (.A(_0759_),
    .B(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__o21bai_1 _5757_ (.A1(_0753_),
    .A2(_0754_),
    .B1_N(_0758_),
    .Y(_0787_));
 sky130_fd_sc_hd__a21oi_1 _5758_ (.A1(_0756_),
    .A2(_0786_),
    .B1(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__nand2_1 _5759_ (.A(_0726_),
    .B(_2986_),
    .Y(_0789_));
 sky130_fd_sc_hd__and4_1 _5760_ (.A(_0726_),
    .B(_0730_),
    .C(_2975_),
    .D(_3030_),
    .X(_0790_));
 sky130_fd_sc_hd__a21o_1 _5761_ (.A1(_0789_),
    .A2(_0753_),
    .B1(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__nor2_1 _5762_ (.A(_0788_),
    .B(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__o21a_1 _5763_ (.A1(_0750_),
    .A2(_0790_),
    .B1(_0749_),
    .X(_0793_));
 sky130_fd_sc_hd__or3_1 _5764_ (.A(_0743_),
    .B(_0746_),
    .C(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__a31o_1 _5765_ (.A1(_0749_),
    .A2(_0752_),
    .A3(_0792_),
    .B1(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__and2_1 _5766_ (.A(_0742_),
    .B(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__a22oi_1 _5767_ (.A1(_0726_),
    .A2(_2711_),
    .B1(_2777_),
    .B2(_0730_),
    .Y(_0797_));
 sky130_fd_sc_hd__nor2_1 _5768_ (.A(_0739_),
    .B(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__o21a_1 _5769_ (.A1(_0740_),
    .A2(_0796_),
    .B1(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__xor2_1 _5770_ (.A(_0737_),
    .B(_0738_),
    .X(_0800_));
 sky130_fd_sc_hd__o21a_1 _5771_ (.A1(_0739_),
    .A2(_0799_),
    .B1(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__o21bai_1 _5772_ (.A1(_0737_),
    .A2(_0738_),
    .B1_N(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__a21oi_1 _5773_ (.A1(_0736_),
    .A2(_0802_),
    .B1(_0734_),
    .Y(_0803_));
 sky130_fd_sc_hd__a22oi_1 _5774_ (.A1(_0727_),
    .A2(_2557_),
    .B1(_2623_),
    .B2(_0731_),
    .Y(_0804_));
 sky130_fd_sc_hd__nor2_1 _5775_ (.A(_0733_),
    .B(_0804_),
    .Y(_0805_));
 sky130_fd_sc_hd__nor2b_1 _5776_ (.A(_0803_),
    .B_N(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__a22oi_1 _5777_ (.A1(_0727_),
    .A2(_2469_),
    .B1(_2568_),
    .B2(_0731_),
    .Y(_0807_));
 sky130_fd_sc_hd__nor2_1 _5778_ (.A(_0732_),
    .B(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__o21a_1 _5779_ (.A1(_0733_),
    .A2(_0806_),
    .B1(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__nand2_1 _5780_ (.A(_0731_),
    .B(_2480_),
    .Y(_0810_));
 sky130_fd_sc_hd__nand2_1 _5781_ (.A(_0727_),
    .B(_3800_),
    .Y(_0811_));
 sky130_fd_sc_hd__xor2_1 _5782_ (.A(_0810_),
    .B(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__o21a_1 _5783_ (.A1(_0732_),
    .A2(_0809_),
    .B1(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__and3_1 _5784_ (.A(_0727_),
    .B(_0731_),
    .C(_3800_),
    .X(_0814_));
 sky130_fd_sc_hd__nor2_1 _5785_ (.A(_0813_),
    .B(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__buf_2 _5786_ (.A(\In2_reg[10] ),
    .X(_0816_));
 sky130_fd_sc_hd__buf_2 _5787_ (.A(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__buf_2 _5788_ (.A(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__buf_2 _5789_ (.A(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__nand4_1 _5790_ (.A(_0819_),
    .B(_3801_),
    .C(_2491_),
    .D(_0722_),
    .Y(_0820_));
 sky130_fd_sc_hd__and3_1 _5791_ (.A(_0819_),
    .B(_3801_),
    .C(_0722_),
    .X(_0821_));
 sky130_fd_sc_hd__a21oi_1 _5792_ (.A1(_3801_),
    .A2(_0722_),
    .B1(_0819_),
    .Y(_0822_));
 sky130_fd_sc_hd__or2_1 _5793_ (.A(_0821_),
    .B(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__nand2_1 _5794_ (.A(_0820_),
    .B(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__a22o_1 _5795_ (.A1(_0819_),
    .A2(_3800_),
    .B1(_2480_),
    .B2(_0722_),
    .X(_0825_));
 sky130_fd_sc_hd__and4_1 _5796_ (.A(_0819_),
    .B(_2568_),
    .C(_2623_),
    .D(_0721_),
    .X(_0826_));
 sky130_fd_sc_hd__and4_1 _5797_ (.A(_0819_),
    .B(_2469_),
    .C(_2568_),
    .D(_0722_),
    .X(_0827_));
 sky130_fd_sc_hd__a22oi_1 _5798_ (.A1(_0819_),
    .A2(_2568_),
    .B1(_2634_),
    .B2(_0722_),
    .Y(_0828_));
 sky130_fd_sc_hd__or2_1 _5799_ (.A(_0826_),
    .B(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__a22oi_1 _5800_ (.A1(_0819_),
    .A2(_2480_),
    .B1(_2568_),
    .B2(_0722_),
    .Y(_0830_));
 sky130_fd_sc_hd__or2_1 _5801_ (.A(_0827_),
    .B(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__and4_1 _5802_ (.A(_2678_),
    .B(_0819_),
    .C(_2623_),
    .D(_0721_),
    .X(_0832_));
 sky130_fd_sc_hd__a22oi_1 _5803_ (.A1(_0819_),
    .A2(_2623_),
    .B1(_0722_),
    .B2(_2678_),
    .Y(_0833_));
 sky130_fd_sc_hd__nor2_1 _5804_ (.A(_0832_),
    .B(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__a22o_1 _5805_ (.A1(_2722_),
    .A2(_0818_),
    .B1(_0721_),
    .B2(_2788_),
    .X(_0835_));
 sky130_fd_sc_hd__and4_1 _5806_ (.A(_2777_),
    .B(_2832_),
    .C(_0818_),
    .D(_0721_),
    .X(_0836_));
 sky130_fd_sc_hd__nand2_1 _5807_ (.A(_2832_),
    .B(_0721_),
    .Y(_0837_));
 sky130_fd_sc_hd__nand2_1 _5808_ (.A(_2865_),
    .B(_0818_),
    .Y(_0838_));
 sky130_fd_sc_hd__nor2_1 _5809_ (.A(_0837_),
    .B(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__a22o_1 _5810_ (.A1(_2832_),
    .A2(_0818_),
    .B1(_0721_),
    .B2(_2865_),
    .X(_0840_));
 sky130_fd_sc_hd__o21ai_1 _5811_ (.A1(_0837_),
    .A2(_0838_),
    .B1(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__a22o_1 _5812_ (.A1(_2909_),
    .A2(_0818_),
    .B1(_0721_),
    .B2(_2997_),
    .X(_0842_));
 sky130_fd_sc_hd__nand2_1 _5813_ (.A(_3041_),
    .B(_0720_),
    .Y(_0843_));
 sky130_fd_sc_hd__nand2_1 _5814_ (.A(_2986_),
    .B(_0817_),
    .Y(_0844_));
 sky130_fd_sc_hd__and4_1 _5815_ (.A(_2986_),
    .B(_3030_),
    .C(_0817_),
    .D(_0720_),
    .X(_0845_));
 sky130_fd_sc_hd__a21o_1 _5816_ (.A1(_0843_),
    .A2(_0844_),
    .B1(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__a22o_1 _5817_ (.A1(_3030_),
    .A2(_0817_),
    .B1(_0720_),
    .B2(_3096_),
    .X(_0847_));
 sky130_fd_sc_hd__nand2_1 _5818_ (.A(_3085_),
    .B(_0817_),
    .Y(_0848_));
 sky130_fd_sc_hd__nand2_1 _5819_ (.A(_3140_),
    .B(_0720_),
    .Y(_0849_));
 sky130_fd_sc_hd__and4_1 _5820_ (.A(_3085_),
    .B(_3129_),
    .C(_0817_),
    .D(_0720_),
    .X(_0850_));
 sky130_fd_sc_hd__a21oi_1 _5821_ (.A1(_0848_),
    .A2(_0849_),
    .B1(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__a22o_1 _5822_ (.A1(_3140_),
    .A2(_0817_),
    .B1(_0720_),
    .B2(_3184_),
    .X(_0852_));
 sky130_fd_sc_hd__and4_1 _5823_ (.A(_3129_),
    .B(_3184_),
    .C(_0817_),
    .D(_0719_),
    .X(_0853_));
 sky130_fd_sc_hd__and3_1 _5824_ (.A(_3162_),
    .B(_3228_),
    .C(_0816_),
    .X(_0854_));
 sky130_fd_sc_hd__a22o_1 _5825_ (.A1(_3173_),
    .A2(_0816_),
    .B1(_0719_),
    .B2(_3228_),
    .X(_0855_));
 sky130_fd_sc_hd__a21bo_1 _5826_ (.A1(_0719_),
    .A2(_0854_),
    .B1_N(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__and4_1 _5827_ (.A(_3228_),
    .B(_3294_),
    .C(_0816_),
    .D(_0719_),
    .X(_0857_));
 sky130_fd_sc_hd__and3_1 _5828_ (.A(_3294_),
    .B(_3349_),
    .C(\M1.U1.U6.u3.instance3_2.Prop_L ),
    .X(_0858_));
 sky130_fd_sc_hd__and3_1 _5829_ (.A(_3349_),
    .B(_3387_),
    .C(_0816_),
    .X(_0859_));
 sky130_fd_sc_hd__a22o_1 _5830_ (.A1(_3349_),
    .A2(_0816_),
    .B1(\M1.U1.U6.u3.instance3_2.Prop_L ),
    .B2(_3387_),
    .X(_0860_));
 sky130_fd_sc_hd__nand2_1 _5831_ (.A(_3380_),
    .B(\In2_reg[10] ),
    .Y(_0861_));
 sky130_fd_sc_hd__nand2_1 _5832_ (.A(_3437_),
    .B(\M1.U1.U6.u3.instance3_2.Prop_L ),
    .Y(_0862_));
 sky130_fd_sc_hd__and4_1 _5833_ (.A(_3380_),
    .B(_3437_),
    .C(\In2_reg[10] ),
    .D(\M1.U1.U6.u3.instance3_2.Prop_L ),
    .X(_0863_));
 sky130_fd_sc_hd__a21o_1 _5834_ (.A1(_0861_),
    .A2(_0862_),
    .B1(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__a22o_1 _5835_ (.A1(_3437_),
    .A2(\In2_reg[10] ),
    .B1(\M1.U1.U6.u3.instance3_2.Prop_L ),
    .B2(_3586_),
    .X(_0865_));
 sky130_fd_sc_hd__o2111a_1 _5836_ (.A1(_3586_),
    .A2(_3536_),
    .B1(\In2_reg[10] ),
    .C1(\M1.U1.U6.u3.instance3_2.Prop_L ),
    .D1(_3503_),
    .X(_0866_));
 sky130_fd_sc_hd__nand2_1 _5837_ (.A(_3596_),
    .B(\In2_reg[10] ),
    .Y(_0867_));
 sky130_fd_sc_hd__o2bb2a_1 _5838_ (.A1_N(_0865_),
    .A2_N(_0866_),
    .B1(_0862_),
    .B2(_0867_),
    .X(_0868_));
 sky130_fd_sc_hd__o21bai_2 _5839_ (.A1(_0864_),
    .A2(_0868_),
    .B1_N(_0863_),
    .Y(_0869_));
 sky130_fd_sc_hd__a22o_1 _5840_ (.A1(_0719_),
    .A2(_0859_),
    .B1(_0860_),
    .B2(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__a22o_1 _5841_ (.A1(_3294_),
    .A2(_0816_),
    .B1(_0719_),
    .B2(_3349_),
    .X(_0871_));
 sky130_fd_sc_hd__a22o_1 _5842_ (.A1(_0816_),
    .A2(_0858_),
    .B1(_0870_),
    .B2(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__a22o_1 _5843_ (.A1(_3228_),
    .A2(_0817_),
    .B1(_0719_),
    .B2(_3294_),
    .X(_0873_));
 sky130_fd_sc_hd__o21a_1 _5844_ (.A1(_0857_),
    .A2(_0872_),
    .B1(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__nor2b_1 _5845_ (.A(_0856_),
    .B_N(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__a21o_1 _5846_ (.A1(_0719_),
    .A2(_0854_),
    .B1(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__or2_1 _5847_ (.A(_0853_),
    .B(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__a31o_1 _5848_ (.A1(_0851_),
    .A2(_0852_),
    .A3(_0877_),
    .B1(_0850_),
    .X(_0878_));
 sky130_fd_sc_hd__o2bb2a_1 _5849_ (.A1_N(_0847_),
    .A2_N(_0878_),
    .B1(_0843_),
    .B2(_0848_),
    .X(_0879_));
 sky130_fd_sc_hd__nor2_1 _5850_ (.A(_0846_),
    .B(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__nand2_1 _5851_ (.A(_2909_),
    .B(_0720_),
    .Y(_0881_));
 sky130_fd_sc_hd__o21bai_1 _5852_ (.A1(_0881_),
    .A2(_0844_),
    .B1_N(_0845_),
    .Y(_0882_));
 sky130_fd_sc_hd__a21oi_1 _5853_ (.A1(_0842_),
    .A2(_0880_),
    .B1(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__and4_1 _5854_ (.A(_2865_),
    .B(_2909_),
    .C(_0818_),
    .D(_0720_),
    .X(_0884_));
 sky130_fd_sc_hd__a21o_1 _5855_ (.A1(_0838_),
    .A2(_0881_),
    .B1(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__o21ba_1 _5856_ (.A1(_0883_),
    .A2(_0885_),
    .B1_N(_0884_),
    .X(_0886_));
 sky130_fd_sc_hd__nor2_1 _5857_ (.A(_0841_),
    .B(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__nand2_1 _5858_ (.A(_2788_),
    .B(_0818_),
    .Y(_0888_));
 sky130_fd_sc_hd__a21oi_1 _5859_ (.A1(_0888_),
    .A2(_0837_),
    .B1(_0836_),
    .Y(_0889_));
 sky130_fd_sc_hd__o21a_1 _5860_ (.A1(_0839_),
    .A2(_0887_),
    .B1(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__or2_1 _5861_ (.A(_0836_),
    .B(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__nand2_1 _5862_ (.A(_2722_),
    .B(_0721_),
    .Y(_0892_));
 sky130_fd_sc_hd__o2bb2a_1 _5863_ (.A1_N(_0835_),
    .A2_N(_0891_),
    .B1(_0892_),
    .B2(_0888_),
    .X(_0893_));
 sky130_fd_sc_hd__nand2_1 _5864_ (.A(_2678_),
    .B(_0818_),
    .Y(_0894_));
 sky130_fd_sc_hd__and4_1 _5865_ (.A(_2678_),
    .B(_2722_),
    .C(_0818_),
    .D(_0721_),
    .X(_0895_));
 sky130_fd_sc_hd__a21o_1 _5866_ (.A1(_0892_),
    .A2(_0894_),
    .B1(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__o21bai_1 _5867_ (.A1(_0893_),
    .A2(_0896_),
    .B1_N(_0895_),
    .Y(_0897_));
 sky130_fd_sc_hd__a21oi_1 _5868_ (.A1(_0834_),
    .A2(_0897_),
    .B1(_0832_),
    .Y(_0898_));
 sky130_fd_sc_hd__or3_1 _5869_ (.A(_0829_),
    .B(_0831_),
    .C(_0898_),
    .X(_0899_));
 sky130_fd_sc_hd__or3b_1 _5870_ (.A(_0826_),
    .B(_0827_),
    .C_N(_0899_),
    .X(_0900_));
 sky130_fd_sc_hd__and3_1 _5871_ (.A(_0820_),
    .B(_0825_),
    .C(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _5872_ (.A0(_0824_),
    .A1(_0823_),
    .S(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__and2b_1 _5873_ (.A_N(_0815_),
    .B(_0902_),
    .X(_0903_));
 sky130_fd_sc_hd__and2b_1 _5874_ (.A_N(_0902_),
    .B(_0815_),
    .X(_0904_));
 sky130_fd_sc_hd__nor2_1 _5875_ (.A(_0903_),
    .B(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__nand2_1 _5876_ (.A(_0731_),
    .B(_0815_),
    .Y(_0906_));
 sky130_fd_sc_hd__a21oi_1 _5877_ (.A1(_0820_),
    .A2(_0825_),
    .B1(_0900_),
    .Y(_0907_));
 sky130_fd_sc_hd__or2_1 _5878_ (.A(_0901_),
    .B(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__a21oi_1 _5879_ (.A1(_0731_),
    .A2(_3800_),
    .B1(_0727_),
    .Y(_0909_));
 sky130_fd_sc_hd__nor2_1 _5880_ (.A(_0814_),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__o21bai_1 _5881_ (.A1(_0810_),
    .A2(_0811_),
    .B1_N(_0813_),
    .Y(_0911_));
 sky130_fd_sc_hd__xnor2_1 _5882_ (.A(_0910_),
    .B(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__o21ba_1 _5883_ (.A1(_0829_),
    .A2(_0898_),
    .B1_N(_0826_),
    .X(_0913_));
 sky130_fd_sc_hd__xnor2_1 _5884_ (.A(_0831_),
    .B(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__or2_1 _5885_ (.A(_0912_),
    .B(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__nor3_1 _5886_ (.A(_0812_),
    .B(_0732_),
    .C(_0809_),
    .Y(_0916_));
 sky130_fd_sc_hd__xnor2_1 _5887_ (.A(_0829_),
    .B(_0898_),
    .Y(_0917_));
 sky130_fd_sc_hd__or3_1 _5888_ (.A(_0813_),
    .B(_0916_),
    .C(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__nor3_1 _5889_ (.A(_0808_),
    .B(_0733_),
    .C(_0806_),
    .Y(_0919_));
 sky130_fd_sc_hd__or2_1 _5890_ (.A(_0809_),
    .B(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__xnor2_1 _5891_ (.A(_0834_),
    .B(_0897_),
    .Y(_0921_));
 sky130_fd_sc_hd__or2_1 _5892_ (.A(_0920_),
    .B(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__and2b_1 _5893_ (.A_N(_0805_),
    .B(_0803_),
    .X(_0923_));
 sky130_fd_sc_hd__or2_1 _5894_ (.A(_0806_),
    .B(_0923_),
    .X(_0924_));
 sky130_fd_sc_hd__xnor2_1 _5895_ (.A(_0893_),
    .B(_0896_),
    .Y(_0925_));
 sky130_fd_sc_hd__nor2_1 _5896_ (.A(_0924_),
    .B(_0925_),
    .Y(_0926_));
 sky130_fd_sc_hd__xnor2_1 _5897_ (.A(_0736_),
    .B(_0802_),
    .Y(_0927_));
 sky130_fd_sc_hd__o21a_1 _5898_ (.A1(_0892_),
    .A2(_0888_),
    .B1(_0835_),
    .X(_0928_));
 sky130_fd_sc_hd__xnor2_1 _5899_ (.A(_0928_),
    .B(_0891_),
    .Y(_0929_));
 sky130_fd_sc_hd__or2_1 _5900_ (.A(_0927_),
    .B(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__nor3_1 _5901_ (.A(_0800_),
    .B(_0739_),
    .C(_0799_),
    .Y(_0931_));
 sky130_fd_sc_hd__nor2_1 _5902_ (.A(_0801_),
    .B(_0931_),
    .Y(_0932_));
 sky130_fd_sc_hd__nor3_1 _5903_ (.A(_0839_),
    .B(_0887_),
    .C(_0889_),
    .Y(_0933_));
 sky130_fd_sc_hd__nor2_1 _5904_ (.A(_0890_),
    .B(_0933_),
    .Y(_0934_));
 sky130_fd_sc_hd__and2_1 _5905_ (.A(_0932_),
    .B(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__nor3_1 _5906_ (.A(_0798_),
    .B(_0740_),
    .C(_0796_),
    .Y(_0936_));
 sky130_fd_sc_hd__or2_1 _5907_ (.A(_0799_),
    .B(_0936_),
    .X(_0937_));
 sky130_fd_sc_hd__xnor2_1 _5908_ (.A(_0841_),
    .B(_0886_),
    .Y(_0938_));
 sky130_fd_sc_hd__or2_1 _5909_ (.A(_0937_),
    .B(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__nor2_1 _5910_ (.A(_0742_),
    .B(_0795_),
    .Y(_0940_));
 sky130_fd_sc_hd__nor2_1 _5911_ (.A(_0796_),
    .B(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__xor2_1 _5912_ (.A(_0883_),
    .B(_0885_),
    .X(_0942_));
 sky130_fd_sc_hd__and2_1 _5913_ (.A(_0941_),
    .B(_0942_),
    .X(_0943_));
 sky130_fd_sc_hd__or2_1 _5914_ (.A(_0790_),
    .B(_0792_),
    .X(_0944_));
 sky130_fd_sc_hd__a21oi_1 _5915_ (.A1(_0752_),
    .A2(_0944_),
    .B1(_0750_),
    .Y(_0945_));
 sky130_fd_sc_hd__o21ba_1 _5916_ (.A1(_0745_),
    .A2(_0945_),
    .B1_N(_0743_),
    .X(_0946_));
 sky130_fd_sc_hd__xnor2_1 _5917_ (.A(_0748_),
    .B(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__o21ai_1 _5918_ (.A1(_0881_),
    .A2(_0844_),
    .B1(_0842_),
    .Y(_0948_));
 sky130_fd_sc_hd__nor2_1 _5919_ (.A(_0845_),
    .B(_0880_),
    .Y(_0949_));
 sky130_fd_sc_hd__xnor2_1 _5920_ (.A(_0948_),
    .B(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__nor2_1 _5921_ (.A(_0947_),
    .B(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__xnor2_1 _5922_ (.A(_0745_),
    .B(_0945_),
    .Y(_0952_));
 sky130_fd_sc_hd__and2_1 _5923_ (.A(_0846_),
    .B(_0879_),
    .X(_0953_));
 sky130_fd_sc_hd__or2_1 _5924_ (.A(_0880_),
    .B(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__or2_1 _5925_ (.A(_0952_),
    .B(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__xnor2_1 _5926_ (.A(_0752_),
    .B(_0944_),
    .Y(_0956_));
 sky130_fd_sc_hd__o21a_1 _5927_ (.A1(_0843_),
    .A2(_0848_),
    .B1(_0847_),
    .X(_0957_));
 sky130_fd_sc_hd__xnor2_1 _5928_ (.A(_0957_),
    .B(_0878_),
    .Y(_0958_));
 sky130_fd_sc_hd__nor2_1 _5929_ (.A(_0956_),
    .B(_0958_),
    .Y(_0959_));
 sky130_fd_sc_hd__and2_1 _5930_ (.A(_0788_),
    .B(_0791_),
    .X(_0960_));
 sky130_fd_sc_hd__or2_1 _5931_ (.A(_0792_),
    .B(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__nand2_1 _5932_ (.A(_0852_),
    .B(_0877_),
    .Y(_0962_));
 sky130_fd_sc_hd__xor2_1 _5933_ (.A(_0851_),
    .B(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__nor2_1 _5934_ (.A(_0961_),
    .B(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__nor2_1 _5935_ (.A(_0758_),
    .B(_0786_),
    .Y(_0965_));
 sky130_fd_sc_hd__xnor2_1 _5936_ (.A(_0756_),
    .B(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__or2b_1 _5937_ (.A(_0853_),
    .B_N(_0852_),
    .X(_0967_));
 sky130_fd_sc_hd__xnor2_1 _5938_ (.A(_0876_),
    .B(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__and2_1 _5939_ (.A(_0966_),
    .B(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__and2_1 _5940_ (.A(_0759_),
    .B(_0785_),
    .X(_0970_));
 sky130_fd_sc_hd__or2_1 _5941_ (.A(_0786_),
    .B(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__xor2_1 _5942_ (.A(_0856_),
    .B(_0874_),
    .X(_0972_));
 sky130_fd_sc_hd__nor2_1 _5943_ (.A(_0971_),
    .B(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__or2_1 _5944_ (.A(_0779_),
    .B(_0781_),
    .X(_0974_));
 sky130_fd_sc_hd__xnor2_1 _5945_ (.A(_0783_),
    .B(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__inv_2 _5946_ (.A(_0873_),
    .Y(_0976_));
 sky130_fd_sc_hd__nor2_1 _5947_ (.A(_0976_),
    .B(_0857_),
    .Y(_0977_));
 sky130_fd_sc_hd__xnor2_1 _5948_ (.A(_0872_),
    .B(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__nor2_1 _5949_ (.A(_0975_),
    .B(_0978_),
    .Y(_0979_));
 sky130_fd_sc_hd__xnor2_1 _5950_ (.A(_0780_),
    .B(_0777_),
    .Y(_0980_));
 sky130_fd_sc_hd__a21bo_1 _5951_ (.A1(_0817_),
    .A2(_0858_),
    .B1_N(_0871_),
    .X(_0981_));
 sky130_fd_sc_hd__xnor2_1 _5952_ (.A(_0870_),
    .B(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__o21ai_1 _5953_ (.A1(_0776_),
    .A2(_0761_),
    .B1(_0760_),
    .Y(_0983_));
 sky130_fd_sc_hd__xnor2_1 _5954_ (.A(_0775_),
    .B(_0983_),
    .Y(_0984_));
 sky130_fd_sc_hd__o21ba_1 _5955_ (.A1(_0860_),
    .A2(_0869_),
    .B1_N(_0870_),
    .X(_0985_));
 sky130_fd_sc_hd__a31oi_2 _5956_ (.A1(_0720_),
    .A2(_0859_),
    .A3(_0869_),
    .B1(_0985_),
    .Y(_0986_));
 sky130_fd_sc_hd__inv_2 _5957_ (.A(_0986_),
    .Y(_0987_));
 sky130_fd_sc_hd__nand2_1 _5958_ (.A(_0984_),
    .B(_0987_),
    .Y(_0988_));
 sky130_fd_sc_hd__xnor2_1 _5959_ (.A(_0764_),
    .B(_0774_),
    .Y(_0989_));
 sky130_fd_sc_hd__xnor2_1 _5960_ (.A(_0864_),
    .B(_0868_),
    .Y(_0990_));
 sky130_fd_sc_hd__nor2_1 _5961_ (.A(_0989_),
    .B(_0990_),
    .Y(_0991_));
 sky130_fd_sc_hd__a21bo_1 _5962_ (.A1(_3393_),
    .A2(_0765_),
    .B1_N(_0766_),
    .X(_0992_));
 sky130_fd_sc_hd__xor2_1 _5963_ (.A(_0992_),
    .B(_0773_),
    .X(_0993_));
 sky130_fd_sc_hd__o21a_1 _5964_ (.A1(_0862_),
    .A2(_0867_),
    .B1(_0865_),
    .X(_0994_));
 sky130_fd_sc_hd__xnor2_1 _5965_ (.A(_0994_),
    .B(_0866_),
    .Y(_0995_));
 sky130_fd_sc_hd__nor2_1 _5966_ (.A(_0993_),
    .B(_0995_),
    .Y(_0996_));
 sky130_fd_sc_hd__and2b_1 _5967_ (.A_N(_0772_),
    .B(_0767_),
    .X(_0997_));
 sky130_fd_sc_hd__xnor2_1 _5968_ (.A(_0997_),
    .B(_0771_),
    .Y(_0998_));
 sky130_fd_sc_hd__nand2_1 _5969_ (.A(_3514_),
    .B(\M1.U1.U6.u3.instance3_2.Prop_L ),
    .Y(_0999_));
 sky130_fd_sc_hd__nand2_1 _5970_ (.A(_3546_),
    .B(_0816_),
    .Y(_1000_));
 sky130_fd_sc_hd__or2_1 _5971_ (.A(_0999_),
    .B(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__and3_1 _5972_ (.A(_3596_),
    .B(_3514_),
    .C(\In2_reg[10] ),
    .X(_1002_));
 sky130_fd_sc_hd__a22o_1 _5973_ (.A1(_0867_),
    .A2(_0999_),
    .B1(_1002_),
    .B2(\M1.U1.U6.u3.instance3_2.Prop_L ),
    .X(_1003_));
 sky130_fd_sc_hd__xnor2_1 _5974_ (.A(_1001_),
    .B(_1003_),
    .Y(_1004_));
 sky130_fd_sc_hd__nor2_1 _5975_ (.A(_0998_),
    .B(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__or2b_1 _5976_ (.A(_0770_),
    .B_N(_0768_),
    .X(_1006_));
 sky130_fd_sc_hd__xnor2_1 _5977_ (.A(_1006_),
    .B(_0769_),
    .Y(_1007_));
 sky130_fd_sc_hd__a22o_1 _5978_ (.A1(_3514_),
    .A2(_0816_),
    .B1(_0719_),
    .B2(_3546_),
    .X(_1008_));
 sky130_fd_sc_hd__and3_1 _5979_ (.A(_1001_),
    .B(_1007_),
    .C(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__nand2_1 _5980_ (.A(_1001_),
    .B(_1008_),
    .Y(_1010_));
 sky130_fd_sc_hd__xor2_1 _5981_ (.A(_1007_),
    .B(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__nand2_1 _5982_ (.A(_0724_),
    .B(_3605_),
    .Y(_1012_));
 sky130_fd_sc_hd__nand2_1 _5983_ (.A(_0728_),
    .B(_3514_),
    .Y(_1013_));
 sky130_fd_sc_hd__a21o_1 _5984_ (.A1(_1012_),
    .A2(_1013_),
    .B1(_0769_),
    .X(_1014_));
 sky130_fd_sc_hd__nand2_1 _5985_ (.A(_0724_),
    .B(_3546_),
    .Y(_1015_));
 sky130_fd_sc_hd__or3_1 _5986_ (.A(_1012_),
    .B(_1013_),
    .C(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__a21o_1 _5987_ (.A1(_1014_),
    .A2(_1016_),
    .B1(_1000_),
    .X(_1017_));
 sky130_fd_sc_hd__nor2_1 _5988_ (.A(_1011_),
    .B(_1017_),
    .Y(_1018_));
 sky130_fd_sc_hd__and2_1 _5989_ (.A(_0998_),
    .B(_1004_),
    .X(_1019_));
 sky130_fd_sc_hd__nor2_1 _5990_ (.A(_1005_),
    .B(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__o21a_1 _5991_ (.A1(_1009_),
    .A2(_1018_),
    .B1(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__and2_1 _5992_ (.A(_0993_),
    .B(_0995_),
    .X(_1022_));
 sky130_fd_sc_hd__nor2_1 _5993_ (.A(_0996_),
    .B(_1022_),
    .Y(_1023_));
 sky130_fd_sc_hd__o21a_1 _5994_ (.A1(_1005_),
    .A2(_1021_),
    .B1(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__and2_1 _5995_ (.A(_0989_),
    .B(_0990_),
    .X(_1025_));
 sky130_fd_sc_hd__nor2_1 _5996_ (.A(_0991_),
    .B(_1025_),
    .Y(_1026_));
 sky130_fd_sc_hd__o21a_1 _5997_ (.A1(_0996_),
    .A2(_1024_),
    .B1(_1026_),
    .X(_1027_));
 sky130_fd_sc_hd__xnor2_1 _5998_ (.A(_0984_),
    .B(_0986_),
    .Y(_1028_));
 sky130_fd_sc_hd__o21ai_1 _5999_ (.A1(_0991_),
    .A2(_1027_),
    .B1(_1028_),
    .Y(_1029_));
 sky130_fd_sc_hd__xnor2_1 _6000_ (.A(_0980_),
    .B(_0982_),
    .Y(_1030_));
 sky130_fd_sc_hd__a21oi_1 _6001_ (.A1(_0988_),
    .A2(_1029_),
    .B1(_1030_),
    .Y(_1031_));
 sky130_fd_sc_hd__a21oi_1 _6002_ (.A1(_0980_),
    .A2(_0982_),
    .B1(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__and2_1 _6003_ (.A(_0975_),
    .B(_0978_),
    .X(_1033_));
 sky130_fd_sc_hd__nor2_1 _6004_ (.A(_0979_),
    .B(_1033_),
    .Y(_1034_));
 sky130_fd_sc_hd__and2b_1 _6005_ (.A_N(_1032_),
    .B(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__and2_1 _6006_ (.A(_0971_),
    .B(_0972_),
    .X(_1036_));
 sky130_fd_sc_hd__nor2_1 _6007_ (.A(_0973_),
    .B(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__o21a_1 _6008_ (.A1(_0979_),
    .A2(_1035_),
    .B1(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__nor2_1 _6009_ (.A(_0966_),
    .B(_0968_),
    .Y(_1039_));
 sky130_fd_sc_hd__nor2_1 _6010_ (.A(_0969_),
    .B(_1039_),
    .Y(_1040_));
 sky130_fd_sc_hd__o21a_1 _6011_ (.A1(_0973_),
    .A2(_1038_),
    .B1(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__and2_1 _6012_ (.A(_0961_),
    .B(_0963_),
    .X(_1042_));
 sky130_fd_sc_hd__or2_1 _6013_ (.A(_0964_),
    .B(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__o21ba_1 _6014_ (.A1(_0969_),
    .A2(_1041_),
    .B1_N(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__and2_1 _6015_ (.A(_0956_),
    .B(_0958_),
    .X(_1045_));
 sky130_fd_sc_hd__nor2_1 _6016_ (.A(_0959_),
    .B(_1045_),
    .Y(_1046_));
 sky130_fd_sc_hd__o21a_1 _6017_ (.A1(_0964_),
    .A2(_1044_),
    .B1(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__nand2_1 _6018_ (.A(_0952_),
    .B(_0954_),
    .Y(_1048_));
 sky130_fd_sc_hd__and2_1 _6019_ (.A(_0955_),
    .B(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__o21ai_1 _6020_ (.A1(_0959_),
    .A2(_1047_),
    .B1(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__and2_1 _6021_ (.A(_0947_),
    .B(_0950_),
    .X(_1051_));
 sky130_fd_sc_hd__or2_1 _6022_ (.A(_0951_),
    .B(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__a21oi_1 _6023_ (.A1(_0955_),
    .A2(_1050_),
    .B1(_1052_),
    .Y(_1053_));
 sky130_fd_sc_hd__nor2_1 _6024_ (.A(_0941_),
    .B(_0942_),
    .Y(_1054_));
 sky130_fd_sc_hd__or2_1 _6025_ (.A(_0943_),
    .B(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__o21ba_1 _6026_ (.A1(_0951_),
    .A2(_1053_),
    .B1_N(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__nand2_1 _6027_ (.A(_0937_),
    .B(_0938_),
    .Y(_1057_));
 sky130_fd_sc_hd__and2_1 _6028_ (.A(_0939_),
    .B(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__o21ai_1 _6029_ (.A1(_0943_),
    .A2(_1056_),
    .B1(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__nor2_1 _6030_ (.A(_0932_),
    .B(_0934_),
    .Y(_1060_));
 sky130_fd_sc_hd__or2_1 _6031_ (.A(_0935_),
    .B(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__a21oi_1 _6032_ (.A1(_0939_),
    .A2(_1059_),
    .B1(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__nand2_1 _6033_ (.A(_0927_),
    .B(_0929_),
    .Y(_1063_));
 sky130_fd_sc_hd__and2_1 _6034_ (.A(_0930_),
    .B(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__o21ai_1 _6035_ (.A1(_0935_),
    .A2(_1062_),
    .B1(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__nand2_1 _6036_ (.A(_0924_),
    .B(_0925_),
    .Y(_1066_));
 sky130_fd_sc_hd__or2b_1 _6037_ (.A(_0926_),
    .B_N(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__a21oi_1 _6038_ (.A1(_0930_),
    .A2(_1065_),
    .B1(_1067_),
    .Y(_1068_));
 sky130_fd_sc_hd__nand2_1 _6039_ (.A(_0920_),
    .B(_0921_),
    .Y(_1069_));
 sky130_fd_sc_hd__and2_1 _6040_ (.A(_0922_),
    .B(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__o21ai_1 _6041_ (.A1(_0926_),
    .A2(_1068_),
    .B1(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__o21ai_1 _6042_ (.A1(_0813_),
    .A2(_0916_),
    .B1(_0917_),
    .Y(_1072_));
 sky130_fd_sc_hd__nand2_1 _6043_ (.A(_0918_),
    .B(_1072_),
    .Y(_1073_));
 sky130_fd_sc_hd__a21o_1 _6044_ (.A1(_0922_),
    .A2(_1071_),
    .B1(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__nand2_1 _6045_ (.A(_0912_),
    .B(_0914_),
    .Y(_1075_));
 sky130_fd_sc_hd__nand2_1 _6046_ (.A(_0915_),
    .B(_1075_),
    .Y(_1076_));
 sky130_fd_sc_hd__a21o_1 _6047_ (.A1(_0918_),
    .A2(_1074_),
    .B1(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__xnor2_1 _6048_ (.A(_0906_),
    .B(_0908_),
    .Y(_1078_));
 sky130_fd_sc_hd__a21oi_1 _6049_ (.A1(_0915_),
    .A2(_1077_),
    .B1(_1078_),
    .Y(_1079_));
 sky130_fd_sc_hd__o21bai_1 _6050_ (.A1(_0906_),
    .A2(_0908_),
    .B1_N(_1079_),
    .Y(_1080_));
 sky130_fd_sc_hd__a21oi_1 _6051_ (.A1(_0905_),
    .A2(_1080_),
    .B1(_0903_),
    .Y(_1081_));
 sky130_fd_sc_hd__nor2_1 _6052_ (.A(_0901_),
    .B(_0821_),
    .Y(_1082_));
 sky130_fd_sc_hd__o21ai_1 _6053_ (.A1(_0723_),
    .A2(_1081_),
    .B1(_1082_),
    .Y(_1083_));
 sky130_fd_sc_hd__xnor2_1 _6054_ (.A(_0564_),
    .B(_0711_),
    .Y(_1084_));
 sky130_fd_sc_hd__xor2_1 _6055_ (.A(_1083_),
    .B(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__nand2_1 _6056_ (.A(_0722_),
    .B(_1082_),
    .Y(_1086_));
 sky130_fd_sc_hd__xor2_1 _6057_ (.A(_1081_),
    .B(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__or3_1 _6058_ (.A(_0571_),
    .B(_0708_),
    .C(_0709_),
    .X(_1088_));
 sky130_fd_sc_hd__and2_1 _6059_ (.A(_0710_),
    .B(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__xnor2_1 _6060_ (.A(_0905_),
    .B(_1080_),
    .Y(_1090_));
 sky130_fd_sc_hd__and3_1 _6061_ (.A(_0707_),
    .B(_0575_),
    .C(_0705_),
    .X(_1091_));
 sky130_fd_sc_hd__or2_1 _6062_ (.A(_0708_),
    .B(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__nor2_1 _6063_ (.A(_1090_),
    .B(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__and3_1 _6064_ (.A(_1078_),
    .B(_0915_),
    .C(_1077_),
    .X(_1094_));
 sky130_fd_sc_hd__or2_1 _6065_ (.A(_1079_),
    .B(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__or2_1 _6066_ (.A(_0577_),
    .B(_0704_),
    .X(_1096_));
 sky130_fd_sc_hd__nand2_1 _6067_ (.A(_0705_),
    .B(_1096_),
    .Y(_1097_));
 sky130_fd_sc_hd__or2_1 _6068_ (.A(_1095_),
    .B(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__nand3_1 _6069_ (.A(_1076_),
    .B(_0918_),
    .C(_1074_),
    .Y(_1099_));
 sky130_fd_sc_hd__nand2_1 _6070_ (.A(_1077_),
    .B(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__nand2_1 _6071_ (.A(_0582_),
    .B(_0583_),
    .Y(_1101_));
 sky130_fd_sc_hd__xnor2_1 _6072_ (.A(_0702_),
    .B(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__nor2_1 _6073_ (.A(_1100_),
    .B(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__nand3_1 _6074_ (.A(_1073_),
    .B(_0922_),
    .C(_1071_),
    .Y(_1104_));
 sky130_fd_sc_hd__nand2_1 _6075_ (.A(_1074_),
    .B(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__xnor2_1 _6076_ (.A(_0584_),
    .B(_0585_),
    .Y(_1106_));
 sky130_fd_sc_hd__xnor2_1 _6077_ (.A(_0700_),
    .B(_1106_),
    .Y(_1107_));
 sky130_fd_sc_hd__nor2_1 _6078_ (.A(_1105_),
    .B(_1107_),
    .Y(_1108_));
 sky130_fd_sc_hd__or3_1 _6079_ (.A(_1070_),
    .B(_0926_),
    .C(_1068_),
    .X(_1109_));
 sky130_fd_sc_hd__and2_1 _6080_ (.A(_1071_),
    .B(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__or3_1 _6081_ (.A(_0698_),
    .B(_0590_),
    .C(_0697_),
    .X(_1111_));
 sky130_fd_sc_hd__and2_1 _6082_ (.A(_0699_),
    .B(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__nand2_1 _6083_ (.A(_1110_),
    .B(_1112_),
    .Y(_1113_));
 sky130_fd_sc_hd__and3_1 _6084_ (.A(_1067_),
    .B(_0930_),
    .C(_1065_),
    .X(_1114_));
 sky130_fd_sc_hd__or2_1 _6085_ (.A(_1068_),
    .B(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__and3_1 _6086_ (.A(_0696_),
    .B(_0595_),
    .C(_0694_),
    .X(_1116_));
 sky130_fd_sc_hd__or2_1 _6087_ (.A(_0697_),
    .B(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__or2_1 _6088_ (.A(_1115_),
    .B(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__or3_1 _6089_ (.A(_1064_),
    .B(_0935_),
    .C(_1062_),
    .X(_1119_));
 sky130_fd_sc_hd__nand2_1 _6090_ (.A(_1065_),
    .B(_1119_),
    .Y(_1120_));
 sky130_fd_sc_hd__or3_1 _6091_ (.A(_0693_),
    .B(_0600_),
    .C(_0691_),
    .X(_1121_));
 sky130_fd_sc_hd__nand2_1 _6092_ (.A(_0694_),
    .B(_1121_),
    .Y(_1122_));
 sky130_fd_sc_hd__nor2_1 _6093_ (.A(_1120_),
    .B(_1122_),
    .Y(_1123_));
 sky130_fd_sc_hd__and3_1 _6094_ (.A(_1061_),
    .B(_0939_),
    .C(_1059_),
    .X(_1124_));
 sky130_fd_sc_hd__or2_1 _6095_ (.A(_1062_),
    .B(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__nor3_1 _6096_ (.A(_0690_),
    .B(_0605_),
    .C(_0688_),
    .Y(_1126_));
 sky130_fd_sc_hd__or3_1 _6097_ (.A(_0691_),
    .B(_1125_),
    .C(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__or3_1 _6098_ (.A(_1058_),
    .B(_0943_),
    .C(_1056_),
    .X(_1128_));
 sky130_fd_sc_hd__nand2_1 _6099_ (.A(_1059_),
    .B(_1128_),
    .Y(_1129_));
 sky130_fd_sc_hd__nor3_1 _6100_ (.A(_0687_),
    .B(_0608_),
    .C(_0685_),
    .Y(_1130_));
 sky130_fd_sc_hd__or2_1 _6101_ (.A(_0688_),
    .B(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__nor2_1 _6102_ (.A(_1129_),
    .B(_1131_),
    .Y(_1132_));
 sky130_fd_sc_hd__or3b_1 _6103_ (.A(_0951_),
    .B(_1053_),
    .C_N(_1055_),
    .X(_1133_));
 sky130_fd_sc_hd__and2b_1 _6104_ (.A_N(_1056_),
    .B(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__xnor2_1 _6105_ (.A(_0684_),
    .B(_0610_),
    .Y(_1135_));
 sky130_fd_sc_hd__nand2_1 _6106_ (.A(_1134_),
    .B(_1135_),
    .Y(_1136_));
 sky130_fd_sc_hd__and3_1 _6107_ (.A(_0955_),
    .B(_1050_),
    .C(_1052_),
    .X(_1137_));
 sky130_fd_sc_hd__nor2_1 _6108_ (.A(_1053_),
    .B(_1137_),
    .Y(_1138_));
 sky130_fd_sc_hd__nor3_1 _6109_ (.A(_0619_),
    .B(_0681_),
    .C(_0682_),
    .Y(_1139_));
 sky130_fd_sc_hd__nor2_1 _6110_ (.A(_0683_),
    .B(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__nand2_1 _6111_ (.A(_1138_),
    .B(_1140_),
    .Y(_1141_));
 sky130_fd_sc_hd__or3_1 _6112_ (.A(_1049_),
    .B(_0959_),
    .C(_1047_),
    .X(_1142_));
 sky130_fd_sc_hd__and2_1 _6113_ (.A(_1050_),
    .B(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__nor3_1 _6114_ (.A(_0680_),
    .B(_0624_),
    .C(_0678_),
    .Y(_1144_));
 sky130_fd_sc_hd__nor2_1 _6115_ (.A(_0681_),
    .B(_1144_),
    .Y(_1145_));
 sky130_fd_sc_hd__nand2_1 _6116_ (.A(_1143_),
    .B(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__nor3_1 _6117_ (.A(_1046_),
    .B(_0964_),
    .C(_1044_),
    .Y(_1147_));
 sky130_fd_sc_hd__nor2_1 _6118_ (.A(_1047_),
    .B(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__nor3_1 _6119_ (.A(_0677_),
    .B(_0628_),
    .C(_0675_),
    .Y(_1149_));
 sky130_fd_sc_hd__nor2_1 _6120_ (.A(_0678_),
    .B(_1149_),
    .Y(_1150_));
 sky130_fd_sc_hd__nand2_1 _6121_ (.A(_1148_),
    .B(_1150_),
    .Y(_1151_));
 sky130_fd_sc_hd__nor2_1 _6122_ (.A(_0969_),
    .B(_1041_),
    .Y(_1152_));
 sky130_fd_sc_hd__xnor2_1 _6123_ (.A(_1043_),
    .B(_1152_),
    .Y(_1153_));
 sky130_fd_sc_hd__nor3_1 _6124_ (.A(_0674_),
    .B(_0633_),
    .C(_0672_),
    .Y(_1154_));
 sky130_fd_sc_hd__or3_1 _6125_ (.A(_0675_),
    .B(_1153_),
    .C(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__nor3_1 _6126_ (.A(_1040_),
    .B(_0973_),
    .C(_1038_),
    .Y(_1156_));
 sky130_fd_sc_hd__or2_1 _6127_ (.A(_1041_),
    .B(_1156_),
    .X(_1157_));
 sky130_fd_sc_hd__nor3_1 _6128_ (.A(_0671_),
    .B(_0637_),
    .C(_0669_),
    .Y(_1158_));
 sky130_fd_sc_hd__or2_1 _6129_ (.A(_0672_),
    .B(_1158_),
    .X(_1159_));
 sky130_fd_sc_hd__nor2_1 _6130_ (.A(_1157_),
    .B(_1159_),
    .Y(_1160_));
 sky130_fd_sc_hd__nor3_1 _6131_ (.A(_1037_),
    .B(_0979_),
    .C(_1035_),
    .Y(_1161_));
 sky130_fd_sc_hd__nor2_1 _6132_ (.A(_1038_),
    .B(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__nor3_1 _6133_ (.A(_0668_),
    .B(_0643_),
    .C(_0666_),
    .Y(_1163_));
 sky130_fd_sc_hd__nor2_1 _6134_ (.A(_0669_),
    .B(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__nand2_1 _6135_ (.A(_1162_),
    .B(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__xnor2_1 _6136_ (.A(_1034_),
    .B(_1032_),
    .Y(_1166_));
 sky130_fd_sc_hd__and3_1 _6137_ (.A(_0665_),
    .B(_0647_),
    .C(_0663_),
    .X(_1167_));
 sky130_fd_sc_hd__or2_1 _6138_ (.A(_0666_),
    .B(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__inv_2 _6139_ (.A(_1168_),
    .Y(_1169_));
 sky130_fd_sc_hd__nand2_1 _6140_ (.A(_1166_),
    .B(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__and3_1 _6141_ (.A(_1030_),
    .B(_0988_),
    .C(_1029_),
    .X(_1171_));
 sky130_fd_sc_hd__or2_1 _6142_ (.A(_1031_),
    .B(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__xnor2_1 _6143_ (.A(_0660_),
    .B(_0662_),
    .Y(_1173_));
 sky130_fd_sc_hd__or2_1 _6144_ (.A(_1172_),
    .B(_1173_),
    .X(_1174_));
 sky130_fd_sc_hd__or3_1 _6145_ (.A(_0991_),
    .B(_1027_),
    .C(_1028_),
    .X(_1175_));
 sky130_fd_sc_hd__nand2_1 _6146_ (.A(_1029_),
    .B(_1175_),
    .Y(_1176_));
 sky130_fd_sc_hd__and2_1 _6147_ (.A(_0656_),
    .B(_0658_),
    .X(_1177_));
 sky130_fd_sc_hd__or2_1 _6148_ (.A(_0659_),
    .B(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__nor2_1 _6149_ (.A(_1176_),
    .B(_1178_),
    .Y(_1179_));
 sky130_fd_sc_hd__nor3_1 _6150_ (.A(_1026_),
    .B(_0996_),
    .C(_1024_),
    .Y(_1180_));
 sky130_fd_sc_hd__nand2_1 _6151_ (.A(_0410_),
    .B(_0655_),
    .Y(_1181_));
 sky130_fd_sc_hd__nand2_1 _6152_ (.A(_0656_),
    .B(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__nor3_1 _6153_ (.A(_1027_),
    .B(_1180_),
    .C(_1182_),
    .Y(_1183_));
 sky130_fd_sc_hd__nor2_1 _6154_ (.A(_1027_),
    .B(_1180_),
    .Y(_1184_));
 sky130_fd_sc_hd__xor2_1 _6155_ (.A(_1184_),
    .B(_1182_),
    .X(_1185_));
 sky130_fd_sc_hd__nor3_1 _6156_ (.A(_1023_),
    .B(_1005_),
    .C(_1021_),
    .Y(_1186_));
 sky130_fd_sc_hd__nor2_1 _6157_ (.A(_1024_),
    .B(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__a22oi_1 _6158_ (.A1(_4142_),
    .A2(_0458_),
    .B1(_0463_),
    .B2(_3556_),
    .Y(_1188_));
 sky130_fd_sc_hd__nor2_1 _6159_ (.A(_0504_),
    .B(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__xnor2_1 _6160_ (.A(_1187_),
    .B(_1189_),
    .Y(_1190_));
 sky130_fd_sc_hd__nand2_1 _6161_ (.A(_4210_),
    .B(_0458_),
    .Y(_1191_));
 sky130_fd_sc_hd__nor3_1 _6162_ (.A(_1020_),
    .B(_1009_),
    .C(_1018_),
    .Y(_1192_));
 sky130_fd_sc_hd__nor2_1 _6163_ (.A(_1021_),
    .B(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__or2b_1 _6164_ (.A(_1191_),
    .B_N(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__nor2_1 _6165_ (.A(_1190_),
    .B(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__a21oi_1 _6166_ (.A1(_1187_),
    .A2(_1189_),
    .B1(_1195_),
    .Y(_1196_));
 sky130_fd_sc_hd__nor2_1 _6167_ (.A(_1185_),
    .B(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__and2_1 _6168_ (.A(_1176_),
    .B(_1178_),
    .X(_1198_));
 sky130_fd_sc_hd__nor2_1 _6169_ (.A(_1179_),
    .B(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__o21a_1 _6170_ (.A1(_1183_),
    .A2(_1197_),
    .B1(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__nand2_1 _6171_ (.A(_1172_),
    .B(_1173_),
    .Y(_1201_));
 sky130_fd_sc_hd__and2_1 _6172_ (.A(_1174_),
    .B(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__o21ai_1 _6173_ (.A1(_1179_),
    .A2(_1200_),
    .B1(_1202_),
    .Y(_1203_));
 sky130_fd_sc_hd__or2_1 _6174_ (.A(_1166_),
    .B(_1169_),
    .X(_1204_));
 sky130_fd_sc_hd__nand2_1 _6175_ (.A(_1170_),
    .B(_1204_),
    .Y(_1205_));
 sky130_fd_sc_hd__a21o_1 _6176_ (.A1(_1174_),
    .A2(_1203_),
    .B1(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__xnor2_1 _6177_ (.A(_1162_),
    .B(_1164_),
    .Y(_1207_));
 sky130_fd_sc_hd__a21o_1 _6178_ (.A1(_1170_),
    .A2(_1206_),
    .B1(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__xor2_1 _6179_ (.A(_1157_),
    .B(_1159_),
    .X(_1209_));
 sky130_fd_sc_hd__a21boi_1 _6180_ (.A1(_1165_),
    .A2(_1208_),
    .B1_N(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__nor2_1 _6181_ (.A(_0675_),
    .B(_1154_),
    .Y(_1211_));
 sky130_fd_sc_hd__xnor2_1 _6182_ (.A(_1153_),
    .B(_1211_),
    .Y(_1212_));
 sky130_fd_sc_hd__o21ai_1 _6183_ (.A1(_1160_),
    .A2(_1210_),
    .B1(_1212_),
    .Y(_1213_));
 sky130_fd_sc_hd__xnor2_1 _6184_ (.A(_1148_),
    .B(_1150_),
    .Y(_1214_));
 sky130_fd_sc_hd__a21o_1 _6185_ (.A1(_1155_),
    .A2(_1213_),
    .B1(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__xnor2_1 _6186_ (.A(_1143_),
    .B(_1145_),
    .Y(_1216_));
 sky130_fd_sc_hd__a21o_1 _6187_ (.A1(_1151_),
    .A2(_1215_),
    .B1(_1216_),
    .X(_1217_));
 sky130_fd_sc_hd__xnor2_1 _6188_ (.A(_1138_),
    .B(_1140_),
    .Y(_1218_));
 sky130_fd_sc_hd__a21o_1 _6189_ (.A1(_1146_),
    .A2(_1217_),
    .B1(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__xnor2_1 _6190_ (.A(_1134_),
    .B(_1135_),
    .Y(_1220_));
 sky130_fd_sc_hd__a21o_1 _6191_ (.A1(_1141_),
    .A2(_1219_),
    .B1(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__xnor2_1 _6192_ (.A(_1129_),
    .B(_1131_),
    .Y(_1222_));
 sky130_fd_sc_hd__a21oi_1 _6193_ (.A1(_1136_),
    .A2(_1221_),
    .B1(_1222_),
    .Y(_1223_));
 sky130_fd_sc_hd__nor2_1 _6194_ (.A(_0691_),
    .B(_1126_),
    .Y(_1224_));
 sky130_fd_sc_hd__xnor2_1 _6195_ (.A(_1125_),
    .B(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__o21ai_1 _6196_ (.A1(_1132_),
    .A2(_1223_),
    .B1(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__xnor2_1 _6197_ (.A(_1120_),
    .B(_1122_),
    .Y(_1227_));
 sky130_fd_sc_hd__a21oi_1 _6198_ (.A1(_1127_),
    .A2(_1226_),
    .B1(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__xor2_1 _6199_ (.A(_1115_),
    .B(_1117_),
    .X(_1229_));
 sky130_fd_sc_hd__o21ai_1 _6200_ (.A1(_1123_),
    .A2(_1228_),
    .B1(_1229_),
    .Y(_1230_));
 sky130_fd_sc_hd__xnor2_1 _6201_ (.A(_1110_),
    .B(_1112_),
    .Y(_1231_));
 sky130_fd_sc_hd__a21o_1 _6202_ (.A1(_1118_),
    .A2(_1230_),
    .B1(_1231_),
    .X(_1232_));
 sky130_fd_sc_hd__xnor2_1 _6203_ (.A(_1105_),
    .B(_1107_),
    .Y(_1233_));
 sky130_fd_sc_hd__a21oi_1 _6204_ (.A1(_1113_),
    .A2(_1232_),
    .B1(_1233_),
    .Y(_1234_));
 sky130_fd_sc_hd__xnor2_1 _6205_ (.A(_1100_),
    .B(_1102_),
    .Y(_1235_));
 sky130_fd_sc_hd__o21ba_1 _6206_ (.A1(_1108_),
    .A2(_1234_),
    .B1_N(_1235_),
    .X(_1236_));
 sky130_fd_sc_hd__xor2_1 _6207_ (.A(_1095_),
    .B(_1097_),
    .X(_1237_));
 sky130_fd_sc_hd__o21ai_1 _6208_ (.A1(_1103_),
    .A2(_1236_),
    .B1(_1237_),
    .Y(_1238_));
 sky130_fd_sc_hd__xnor2_1 _6209_ (.A(_1090_),
    .B(_1092_),
    .Y(_1239_));
 sky130_fd_sc_hd__a21oi_1 _6210_ (.A1(_1098_),
    .A2(_1238_),
    .B1(_1239_),
    .Y(_1240_));
 sky130_fd_sc_hd__xor2_1 _6211_ (.A(_1087_),
    .B(_1089_),
    .X(_1241_));
 sky130_fd_sc_hd__o21a_1 _6212_ (.A1(_1093_),
    .A2(_1240_),
    .B1(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__a21oi_1 _6213_ (.A1(_1087_),
    .A2(_1089_),
    .B1(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__and2b_1 _6214_ (.A_N(_1084_),
    .B(_1083_),
    .X(_1244_));
 sky130_fd_sc_hd__o21ba_1 _6215_ (.A1(_1085_),
    .A2(_1243_),
    .B1_N(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__xnor2_1 _6216_ (.A(_0712_),
    .B(_0554_),
    .Y(_1246_));
 sky130_fd_sc_hd__and2b_1 _6217_ (.A_N(_1245_),
    .B(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__nor3_1 _6218_ (.A(_0552_),
    .B(_0713_),
    .C(_0715_),
    .Y(_1248_));
 sky130_fd_sc_hd__nor2_1 _6219_ (.A(_0716_),
    .B(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__and2_1 _6220_ (.A(_1247_),
    .B(_1249_),
    .X(_1250_));
 sky130_fd_sc_hd__buf_2 _6221_ (.A(\M1.U1.U4.u2.instance15_14.Prop_L ),
    .X(_1251_));
 sky130_fd_sc_hd__clkbuf_2 _6222_ (.A(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__buf_2 _6223_ (.A(_1252_),
    .X(_1253_));
 sky130_fd_sc_hd__buf_2 _6224_ (.A(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__buf_2 _6225_ (.A(\In2_reg[6] ),
    .X(_1255_));
 sky130_fd_sc_hd__buf_2 _6226_ (.A(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__buf_2 _6227_ (.A(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__buf_2 _6228_ (.A(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__and3_1 _6229_ (.A(_1254_),
    .B(_3801_),
    .C(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__a21oi_1 _6230_ (.A1(_1254_),
    .A2(_3801_),
    .B1(_1258_),
    .Y(_1260_));
 sky130_fd_sc_hd__or2_1 _6231_ (.A(_1259_),
    .B(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__nand2_1 _6232_ (.A(_1254_),
    .B(_2480_),
    .Y(_1262_));
 sky130_fd_sc_hd__nand2_1 _6233_ (.A(_1258_),
    .B(_2568_),
    .Y(_1263_));
 sky130_fd_sc_hd__nand2_1 _6234_ (.A(_1254_),
    .B(_2623_),
    .Y(_1264_));
 sky130_fd_sc_hd__and4_1 _6235_ (.A(_2678_),
    .B(_1254_),
    .C(_1258_),
    .D(_2623_),
    .X(_1265_));
 sky130_fd_sc_hd__and4_1 _6236_ (.A(_2667_),
    .B(_2722_),
    .C(_1254_),
    .D(_1258_),
    .X(_1266_));
 sky130_fd_sc_hd__nand2_1 _6237_ (.A(_2722_),
    .B(_1253_),
    .Y(_1267_));
 sky130_fd_sc_hd__a21boi_1 _6238_ (.A1(_2678_),
    .A2(_1258_),
    .B1_N(_1267_),
    .Y(_1268_));
 sky130_fd_sc_hd__or2_1 _6239_ (.A(_1266_),
    .B(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__a22o_1 _6240_ (.A1(_2788_),
    .A2(_1254_),
    .B1(_1258_),
    .B2(_2722_),
    .X(_1270_));
 sky130_fd_sc_hd__nand2_1 _6241_ (.A(_2832_),
    .B(_1253_),
    .Y(_1271_));
 sky130_fd_sc_hd__nand2_1 _6242_ (.A(_2788_),
    .B(_1257_),
    .Y(_1272_));
 sky130_fd_sc_hd__and4_1 _6243_ (.A(_2788_),
    .B(_2832_),
    .C(_1253_),
    .D(_1257_),
    .X(_1273_));
 sky130_fd_sc_hd__a21o_1 _6244_ (.A1(_1271_),
    .A2(_1272_),
    .B1(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__a22o_1 _6245_ (.A1(_2865_),
    .A2(_1253_),
    .B1(_1257_),
    .B2(_2832_),
    .X(_1275_));
 sky130_fd_sc_hd__and3_1 _6246_ (.A(_2854_),
    .B(_2898_),
    .C(_1253_),
    .X(_1276_));
 sky130_fd_sc_hd__nand2_1 _6247_ (.A(_2854_),
    .B(_1257_),
    .Y(_1277_));
 sky130_fd_sc_hd__nand2_1 _6248_ (.A(_2909_),
    .B(_1253_),
    .Y(_1278_));
 sky130_fd_sc_hd__a22o_1 _6249_ (.A1(_1277_),
    .A2(_1278_),
    .B1(_1276_),
    .B2(_1257_),
    .X(_1279_));
 sky130_fd_sc_hd__and4_1 _6250_ (.A(_2909_),
    .B(_2986_),
    .C(_1253_),
    .D(_1257_),
    .X(_1280_));
 sky130_fd_sc_hd__and4_1 _6251_ (.A(_2975_),
    .B(_3030_),
    .C(_1252_),
    .D(_1256_),
    .X(_1281_));
 sky130_fd_sc_hd__a22oi_1 _6252_ (.A1(_3030_),
    .A2(_1253_),
    .B1(_1257_),
    .B2(_2986_),
    .Y(_1282_));
 sky130_fd_sc_hd__nor2_1 _6253_ (.A(_1281_),
    .B(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__and4_1 _6254_ (.A(_3019_),
    .B(_3085_),
    .C(_1252_),
    .D(_1256_),
    .X(_1284_));
 sky130_fd_sc_hd__nand4_1 _6255_ (.A(_3074_),
    .B(_3129_),
    .C(_1252_),
    .D(_1256_),
    .Y(_1285_));
 sky130_fd_sc_hd__a22o_1 _6256_ (.A1(_3173_),
    .A2(_1252_),
    .B1(_1256_),
    .B2(_3118_),
    .X(_1286_));
 sky130_fd_sc_hd__nand2_1 _6257_ (.A(_3173_),
    .B(_1256_),
    .Y(_1287_));
 sky130_fd_sc_hd__nand2_1 _6258_ (.A(_3228_),
    .B(_1252_),
    .Y(_1288_));
 sky130_fd_sc_hd__and4_1 _6259_ (.A(_3162_),
    .B(_3217_),
    .C(_1252_),
    .D(_1255_),
    .X(_1289_));
 sky130_fd_sc_hd__a21o_1 _6260_ (.A1(_1287_),
    .A2(_1288_),
    .B1(_1289_),
    .X(_1290_));
 sky130_fd_sc_hd__a22o_1 _6261_ (.A1(_3294_),
    .A2(_1251_),
    .B1(_1256_),
    .B2(_3217_),
    .X(_1291_));
 sky130_fd_sc_hd__nand2_1 _6262_ (.A(_3338_),
    .B(_1251_),
    .Y(_1292_));
 sky130_fd_sc_hd__nand2_1 _6263_ (.A(_3380_),
    .B(\In2_reg[6] ),
    .Y(_1293_));
 sky130_fd_sc_hd__and4_1 _6264_ (.A(\In1_reg[4] ),
    .B(_3426_),
    .C(\M1.U1.U4.u2.instance15_14.Prop_L ),
    .D(\In2_reg[6] ),
    .X(_1294_));
 sky130_fd_sc_hd__and4_1 _6265_ (.A(_3437_),
    .B(_3586_),
    .C(_1251_),
    .D(\In2_reg[6] ),
    .X(_1295_));
 sky130_fd_sc_hd__nand4_1 _6266_ (.A(_3437_),
    .B(_3576_),
    .C(\M1.U1.U4.u2.instance15_14.Prop_L ),
    .D(\In2_reg[6] ),
    .Y(_1296_));
 sky130_fd_sc_hd__a22o_1 _6267_ (.A1(_3576_),
    .A2(\M1.U1.U4.u2.instance15_14.Prop_L ),
    .B1(\In2_reg[6] ),
    .B2(_3426_),
    .X(_1297_));
 sky130_fd_sc_hd__o2111a_1 _6268_ (.A1(_3576_),
    .A2(_3536_),
    .B1(\M1.U1.U4.u2.instance15_14.Prop_L ),
    .C1(\In2_reg[6] ),
    .D1(net126),
    .X(_1298_));
 sky130_fd_sc_hd__and3_1 _6269_ (.A(_1296_),
    .B(_1297_),
    .C(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__nand2_1 _6270_ (.A(_3437_),
    .B(\M1.U1.U4.u2.instance15_14.Prop_L ),
    .Y(_1300_));
 sky130_fd_sc_hd__a21o_1 _6271_ (.A1(_1293_),
    .A2(_1300_),
    .B1(_1294_),
    .X(_1301_));
 sky130_fd_sc_hd__o21ba_1 _6272_ (.A1(_1295_),
    .A2(_1299_),
    .B1_N(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__or2_1 _6273_ (.A(_1292_),
    .B(_1293_),
    .X(_1303_));
 sky130_fd_sc_hd__a22o_1 _6274_ (.A1(_3380_),
    .A2(_1251_),
    .B1(_1255_),
    .B2(_3338_),
    .X(_1304_));
 sky130_fd_sc_hd__o211a_1 _6275_ (.A1(_1294_),
    .A2(_1302_),
    .B1(_1303_),
    .C1(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__o21ba_1 _6276_ (.A1(_1292_),
    .A2(_1293_),
    .B1_N(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__nand2_1 _6277_ (.A(_3294_),
    .B(_1255_),
    .Y(_1307_));
 sky130_fd_sc_hd__and4_1 _6278_ (.A(_3283_),
    .B(_3349_),
    .C(_1251_),
    .D(_1255_),
    .X(_1308_));
 sky130_fd_sc_hd__a21o_1 _6279_ (.A1(_1307_),
    .A2(_1292_),
    .B1(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__o21bai_1 _6280_ (.A1(_1306_),
    .A2(_1309_),
    .B1_N(_1308_),
    .Y(_1310_));
 sky130_fd_sc_hd__o2bb2a_1 _6281_ (.A1_N(_1291_),
    .A2_N(_1310_),
    .B1(_1288_),
    .B2(_1307_),
    .X(_1311_));
 sky130_fd_sc_hd__nor2_1 _6282_ (.A(_1290_),
    .B(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__nand2_1 _6283_ (.A(_3118_),
    .B(_1252_),
    .Y(_1313_));
 sky130_fd_sc_hd__nor2_1 _6284_ (.A(_1313_),
    .B(_1287_),
    .Y(_1314_));
 sky130_fd_sc_hd__a211o_1 _6285_ (.A1(_1286_),
    .A2(_1312_),
    .B1(_1314_),
    .C1(_1289_),
    .X(_1315_));
 sky130_fd_sc_hd__a22o_1 _6286_ (.A1(_3129_),
    .A2(_1252_),
    .B1(_1256_),
    .B2(_3074_),
    .X(_1316_));
 sky130_fd_sc_hd__nand3_1 _6287_ (.A(_1285_),
    .B(_1315_),
    .C(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__nand2_1 _6288_ (.A(_1285_),
    .B(_1317_),
    .Y(_1318_));
 sky130_fd_sc_hd__a22oi_1 _6289_ (.A1(_3085_),
    .A2(_1252_),
    .B1(_1256_),
    .B2(_3030_),
    .Y(_1319_));
 sky130_fd_sc_hd__o21ba_1 _6290_ (.A1(_1284_),
    .A2(_1318_),
    .B1_N(_1319_),
    .X(_1320_));
 sky130_fd_sc_hd__a21o_1 _6291_ (.A1(_1283_),
    .A2(_1320_),
    .B1(_1281_),
    .X(_1321_));
 sky130_fd_sc_hd__a22o_1 _6292_ (.A1(_2986_),
    .A2(_1253_),
    .B1(_1257_),
    .B2(_2909_),
    .X(_1322_));
 sky130_fd_sc_hd__o21a_1 _6293_ (.A1(_1280_),
    .A2(_1321_),
    .B1(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__nor2b_1 _6294_ (.A(_1279_),
    .B_N(_1323_),
    .Y(_1324_));
 sky130_fd_sc_hd__a21o_1 _6295_ (.A1(_1257_),
    .A2(_1276_),
    .B1(_1324_),
    .X(_1325_));
 sky130_fd_sc_hd__o2bb2a_1 _6296_ (.A1_N(_1275_),
    .A2_N(_1325_),
    .B1(_1271_),
    .B2(_1277_),
    .X(_1326_));
 sky130_fd_sc_hd__nor2_1 _6297_ (.A(_1274_),
    .B(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__nor2_1 _6298_ (.A(_1267_),
    .B(_1272_),
    .Y(_1328_));
 sky130_fd_sc_hd__a211o_1 _6299_ (.A1(_1270_),
    .A2(_1327_),
    .B1(_1328_),
    .C1(_1273_),
    .X(_1329_));
 sky130_fd_sc_hd__nor2b_1 _6300_ (.A(_1269_),
    .B_N(_1329_),
    .Y(_1330_));
 sky130_fd_sc_hd__a22oi_1 _6301_ (.A1(_2678_),
    .A2(_1254_),
    .B1(_1258_),
    .B2(_2623_),
    .Y(_1331_));
 sky130_fd_sc_hd__or2_1 _6302_ (.A(_1265_),
    .B(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__o21ba_1 _6303_ (.A1(_1266_),
    .A2(_1330_),
    .B1_N(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__nand2_1 _6304_ (.A(_1263_),
    .B(_1264_),
    .Y(_1334_));
 sky130_fd_sc_hd__or2_1 _6305_ (.A(_1263_),
    .B(_1264_),
    .X(_1335_));
 sky130_fd_sc_hd__o211a_1 _6306_ (.A1(_1265_),
    .A2(_1333_),
    .B1(_1334_),
    .C1(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__o21ba_1 _6307_ (.A1(_1263_),
    .A2(_1264_),
    .B1_N(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__a22o_1 _6308_ (.A1(_1258_),
    .A2(_2480_),
    .B1(_2579_),
    .B2(_1254_),
    .X(_1338_));
 sky130_fd_sc_hd__o21ai_1 _6309_ (.A1(_1262_),
    .A2(_1263_),
    .B1(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__o22ai_2 _6310_ (.A1(_1262_),
    .A2(_1263_),
    .B1(_1337_),
    .B2(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__nand2_1 _6311_ (.A(_3800_),
    .B(_1258_),
    .Y(_1341_));
 sky130_fd_sc_hd__nand2_1 _6312_ (.A(_1341_),
    .B(_1262_),
    .Y(_1342_));
 sky130_fd_sc_hd__nor2_1 _6313_ (.A(_1341_),
    .B(_1262_),
    .Y(_1343_));
 sky130_fd_sc_hd__a21oi_1 _6314_ (.A1(_1340_),
    .A2(_1342_),
    .B1(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__o21ba_1 _6315_ (.A1(_1261_),
    .A2(_1344_),
    .B1_N(_1259_),
    .X(_1345_));
 sky130_fd_sc_hd__and2_1 _6316_ (.A(_1254_),
    .B(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__clkbuf_2 _6317_ (.A(\M1.U1.U3.u2.instance13_12.Prop_L ),
    .X(_1347_));
 sky130_fd_sc_hd__buf_2 _6318_ (.A(_1347_),
    .X(_1348_));
 sky130_fd_sc_hd__clkbuf_2 _6319_ (.A(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__buf_2 _6320_ (.A(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__xor2_1 _6321_ (.A(_1261_),
    .B(_1344_),
    .X(_1351_));
 sky130_fd_sc_hd__buf_6 _6322_ (.A(\In2_reg[4] ),
    .X(_1352_));
 sky130_fd_sc_hd__buf_2 _6323_ (.A(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__clkbuf_2 _6324_ (.A(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__buf_2 _6325_ (.A(_1354_),
    .X(_1355_));
 sky130_fd_sc_hd__nand2_1 _6326_ (.A(_3800_),
    .B(_1355_),
    .Y(_1356_));
 sky130_fd_sc_hd__nand2_1 _6327_ (.A(_3800_),
    .B(_1350_),
    .Y(_1357_));
 sky130_fd_sc_hd__xor2_1 _6328_ (.A(_1355_),
    .B(_1357_),
    .X(_1358_));
 sky130_fd_sc_hd__nand2_1 _6329_ (.A(_2480_),
    .B(_1350_),
    .Y(_1359_));
 sky130_fd_sc_hd__nand2_1 _6330_ (.A(_1356_),
    .B(_1359_),
    .Y(_1360_));
 sky130_fd_sc_hd__nand2_1 _6331_ (.A(_2557_),
    .B(_1355_),
    .Y(_1361_));
 sky130_fd_sc_hd__a22o_1 _6332_ (.A1(_2568_),
    .A2(_1350_),
    .B1(_1355_),
    .B2(_2469_),
    .X(_1362_));
 sky130_fd_sc_hd__nand2_1 _6333_ (.A(_2612_),
    .B(_1350_),
    .Y(_1363_));
 sky130_fd_sc_hd__xor2_1 _6334_ (.A(_1361_),
    .B(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__a22o_1 _6335_ (.A1(_2667_),
    .A2(_1350_),
    .B1(_1355_),
    .B2(_2612_),
    .X(_1365_));
 sky130_fd_sc_hd__nand2_1 _6336_ (.A(_2711_),
    .B(_1350_),
    .Y(_1366_));
 sky130_fd_sc_hd__nand2_1 _6337_ (.A(_2667_),
    .B(_1355_),
    .Y(_1367_));
 sky130_fd_sc_hd__and4_1 _6338_ (.A(_2667_),
    .B(_2711_),
    .C(_1350_),
    .D(_1355_),
    .X(_1368_));
 sky130_fd_sc_hd__a21o_1 _6339_ (.A1(_1366_),
    .A2(_1367_),
    .B1(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__a22o_1 _6340_ (.A1(_2788_),
    .A2(_1349_),
    .B1(_1355_),
    .B2(_2711_),
    .X(_1370_));
 sky130_fd_sc_hd__nand2_1 _6341_ (.A(_2777_),
    .B(_1355_),
    .Y(_1371_));
 sky130_fd_sc_hd__nand2_1 _6342_ (.A(_2821_),
    .B(_1349_),
    .Y(_1372_));
 sky130_fd_sc_hd__and4_1 _6343_ (.A(_2777_),
    .B(_2821_),
    .C(_1349_),
    .D(_1355_),
    .X(_1373_));
 sky130_fd_sc_hd__a21o_1 _6344_ (.A1(_1371_),
    .A2(_1372_),
    .B1(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__and4_1 _6345_ (.A(_2821_),
    .B(_2865_),
    .C(_1349_),
    .D(_1354_),
    .X(_1375_));
 sky130_fd_sc_hd__and3_1 _6346_ (.A(_2854_),
    .B(_2909_),
    .C(_1354_),
    .X(_1376_));
 sky130_fd_sc_hd__a22o_1 _6347_ (.A1(_2909_),
    .A2(_1349_),
    .B1(_1354_),
    .B2(_2854_),
    .X(_1377_));
 sky130_fd_sc_hd__and4_1 _6348_ (.A(_2898_),
    .B(_2975_),
    .C(_1349_),
    .D(_1354_),
    .X(_1378_));
 sky130_fd_sc_hd__and2_1 _6349_ (.A(_2975_),
    .B(_1348_),
    .X(_1379_));
 sky130_fd_sc_hd__and2_1 _6350_ (.A(_3019_),
    .B(_1354_),
    .X(_1380_));
 sky130_fd_sc_hd__a21o_1 _6351_ (.A1(_3085_),
    .A2(_1348_),
    .B1(_1380_),
    .X(_1381_));
 sky130_fd_sc_hd__nand2_1 _6352_ (.A(_3118_),
    .B(_1348_),
    .Y(_1382_));
 sky130_fd_sc_hd__nand2_1 _6353_ (.A(_3074_),
    .B(_1354_),
    .Y(_1383_));
 sky130_fd_sc_hd__and4_1 _6354_ (.A(_3074_),
    .B(_3118_),
    .C(_1348_),
    .D(_1353_),
    .X(_1384_));
 sky130_fd_sc_hd__a21o_1 _6355_ (.A1(_1382_),
    .A2(_1383_),
    .B1(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__a22o_1 _6356_ (.A1(_3173_),
    .A2(_1348_),
    .B1(_1353_),
    .B2(_3118_),
    .X(_1386_));
 sky130_fd_sc_hd__nand2_1 _6357_ (.A(_3217_),
    .B(_1347_),
    .Y(_1387_));
 sky130_fd_sc_hd__nand2_1 _6358_ (.A(_3283_),
    .B(_1353_),
    .Y(_1388_));
 sky130_fd_sc_hd__and4_1 _6359_ (.A(_3283_),
    .B(_3338_),
    .C(_1347_),
    .D(_1352_),
    .X(_1389_));
 sky130_fd_sc_hd__and4_1 _6360_ (.A(_3338_),
    .B(_3380_),
    .C(_1347_),
    .D(_1353_),
    .X(_1390_));
 sky130_fd_sc_hd__and4_1 _6361_ (.A(\In1_reg[4] ),
    .B(_3426_),
    .C(\M1.U1.U3.u2.instance13_12.Prop_L ),
    .D(_1352_),
    .X(_1391_));
 sky130_fd_sc_hd__inv_2 _6362_ (.A(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__a22o_1 _6363_ (.A1(_3437_),
    .A2(_1347_),
    .B1(_1352_),
    .B2(_3380_),
    .X(_1393_));
 sky130_fd_sc_hd__and4_1 _6364_ (.A(\In1_reg[1] ),
    .B(_3536_),
    .C(\M1.U1.U3.u2.instance13_12.Prop_L ),
    .D(\In2_reg[4] ),
    .X(_1394_));
 sky130_fd_sc_hd__and4_1 _6365_ (.A(\In1_reg[2] ),
    .B(\In1_reg[1] ),
    .C(\M1.U1.U3.u2.instance13_12.Prop_L ),
    .D(_1352_),
    .X(_1395_));
 sky130_fd_sc_hd__and4_1 _6366_ (.A(\In1_reg[3] ),
    .B(_3576_),
    .C(\M1.U1.U3.u2.instance13_12.Prop_L ),
    .D(_1352_),
    .X(_1396_));
 sky130_fd_sc_hd__a211o_1 _6367_ (.A1(_3426_),
    .A2(_1394_),
    .B1(_1395_),
    .C1(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__and3_1 _6368_ (.A(_1392_),
    .B(_1393_),
    .C(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__nand4_1 _6369_ (.A(_3338_),
    .B(_3380_),
    .C(_1347_),
    .D(_1353_),
    .Y(_1399_));
 sky130_fd_sc_hd__a22o_1 _6370_ (.A1(_3380_),
    .A2(_1347_),
    .B1(_1352_),
    .B2(_3338_),
    .X(_1400_));
 sky130_fd_sc_hd__o211a_1 _6371_ (.A1(_1391_),
    .A2(_1398_),
    .B1(_1399_),
    .C1(_1400_),
    .X(_1401_));
 sky130_fd_sc_hd__nand2_1 _6372_ (.A(_3338_),
    .B(_1347_),
    .Y(_1402_));
 sky130_fd_sc_hd__a21o_1 _6373_ (.A1(_1388_),
    .A2(_1402_),
    .B1(_1389_),
    .X(_1403_));
 sky130_fd_sc_hd__o21ba_1 _6374_ (.A1(_1390_),
    .A2(_1401_),
    .B1_N(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__or2_1 _6375_ (.A(_1387_),
    .B(_1388_),
    .X(_1405_));
 sky130_fd_sc_hd__a22o_1 _6376_ (.A1(_3283_),
    .A2(_1347_),
    .B1(_1353_),
    .B2(_3217_),
    .X(_1406_));
 sky130_fd_sc_hd__o211a_1 _6377_ (.A1(_1389_),
    .A2(_1404_),
    .B1(_1405_),
    .C1(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__o21ba_2 _6378_ (.A1(_1387_),
    .A2(_1388_),
    .B1_N(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__nand2_1 _6379_ (.A(_3162_),
    .B(_1353_),
    .Y(_1409_));
 sky130_fd_sc_hd__and4_1 _6380_ (.A(_3162_),
    .B(_3217_),
    .C(_1348_),
    .D(_1353_),
    .X(_1410_));
 sky130_fd_sc_hd__a21o_1 _6381_ (.A1(_1409_),
    .A2(_1387_),
    .B1(_1410_),
    .X(_1411_));
 sky130_fd_sc_hd__o21bai_4 _6382_ (.A1(_1411_),
    .A2(_1408_),
    .B1_N(_1410_),
    .Y(_1412_));
 sky130_fd_sc_hd__o2bb2a_4 _6383_ (.A1_N(_1386_),
    .A2_N(_1412_),
    .B1(_1382_),
    .B2(_1409_),
    .X(_1413_));
 sky130_fd_sc_hd__nor2_1 _6384_ (.A(_1385_),
    .B(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__and3_1 _6385_ (.A(_3074_),
    .B(_1348_),
    .C(_1380_),
    .X(_1415_));
 sky130_fd_sc_hd__a211o_1 _6386_ (.A1(_1381_),
    .A2(_1414_),
    .B1(_1415_),
    .C1(_1384_),
    .X(_1416_));
 sky130_fd_sc_hd__a22o_1 _6387_ (.A1(_3030_),
    .A2(_1348_),
    .B1(_1354_),
    .B2(_2975_),
    .X(_1417_));
 sky130_fd_sc_hd__a22o_1 _6388_ (.A1(_1379_),
    .A2(_1380_),
    .B1(_1416_),
    .B2(_1417_),
    .X(_1418_));
 sky130_fd_sc_hd__a21o_1 _6389_ (.A1(_2898_),
    .A2(_1354_),
    .B1(_1379_),
    .X(_1419_));
 sky130_fd_sc_hd__o21a_1 _6390_ (.A1(_1378_),
    .A2(_1418_),
    .B1(_1419_),
    .X(_1420_));
 sky130_fd_sc_hd__a22o_1 _6391_ (.A1(_1349_),
    .A2(_1376_),
    .B1(_1377_),
    .B2(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__a22o_1 _6392_ (.A1(_2865_),
    .A2(_1349_),
    .B1(_1354_),
    .B2(_2821_),
    .X(_1422_));
 sky130_fd_sc_hd__o21ai_2 _6393_ (.A1(_1375_),
    .A2(_1421_),
    .B1(_1422_),
    .Y(_1423_));
 sky130_fd_sc_hd__o21bai_1 _6394_ (.A1(_1423_),
    .A2(_1374_),
    .B1_N(_1373_),
    .Y(_1424_));
 sky130_fd_sc_hd__o2bb2a_2 _6395_ (.A1_N(_1370_),
    .A2_N(_1424_),
    .B1(_1366_),
    .B2(_1371_),
    .X(_1425_));
 sky130_fd_sc_hd__nor2_1 _6396_ (.A(_1369_),
    .B(_1425_),
    .Y(_1426_));
 sky130_fd_sc_hd__nor2_1 _6397_ (.A(_1363_),
    .B(_1367_),
    .Y(_1427_));
 sky130_fd_sc_hd__a211o_1 _6398_ (.A1(_1365_),
    .A2(_1426_),
    .B1(_1427_),
    .C1(_1368_),
    .X(_1428_));
 sky130_fd_sc_hd__a2bb2o_1 _6399_ (.A1_N(_1361_),
    .A2_N(_1363_),
    .B1(_1364_),
    .B2(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__a2bb2o_2 _6400_ (.A1_N(_1359_),
    .A2_N(_1361_),
    .B1(_1362_),
    .B2(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__nor2_1 _6401_ (.A(_1356_),
    .B(_1359_),
    .Y(_1431_));
 sky130_fd_sc_hd__a21oi_2 _6402_ (.A1(_1360_),
    .A2(_1430_),
    .B1(_1431_),
    .Y(_1432_));
 sky130_fd_sc_hd__or2_1 _6403_ (.A(_1358_),
    .B(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__nand2_1 _6404_ (.A(_1356_),
    .B(_1433_),
    .Y(_1434_));
 sky130_fd_sc_hd__and3_1 _6405_ (.A(_1350_),
    .B(_1356_),
    .C(_1433_),
    .X(_1435_));
 sky130_fd_sc_hd__or2b_1 _6406_ (.A(_1343_),
    .B_N(_1342_),
    .X(_1436_));
 sky130_fd_sc_hd__xnor2_1 _6407_ (.A(_1340_),
    .B(_1436_),
    .Y(_1437_));
 sky130_fd_sc_hd__and2_1 _6408_ (.A(_1435_),
    .B(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__nand2_1 _6409_ (.A(_1358_),
    .B(_1432_),
    .Y(_1439_));
 sky130_fd_sc_hd__and2_1 _6410_ (.A(_1433_),
    .B(_1439_),
    .X(_1440_));
 sky130_fd_sc_hd__xor2_1 _6411_ (.A(_1337_),
    .B(_1339_),
    .X(_1441_));
 sky130_fd_sc_hd__and2_1 _6412_ (.A(_1440_),
    .B(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__or2b_1 _6413_ (.A(_1431_),
    .B_N(_1360_),
    .X(_1443_));
 sky130_fd_sc_hd__xnor2_1 _6414_ (.A(_1443_),
    .B(_1430_),
    .Y(_1444_));
 sky130_fd_sc_hd__a211oi_1 _6415_ (.A1(_1335_),
    .A2(_1334_),
    .B1(_1333_),
    .C1(_1265_),
    .Y(_1445_));
 sky130_fd_sc_hd__nor2_1 _6416_ (.A(_1336_),
    .B(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__and2_1 _6417_ (.A(_1444_),
    .B(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__o21ai_1 _6418_ (.A1(_1359_),
    .A2(_1361_),
    .B1(_1362_),
    .Y(_1448_));
 sky130_fd_sc_hd__xnor2_1 _6419_ (.A(_1448_),
    .B(_1429_),
    .Y(_1449_));
 sky130_fd_sc_hd__or2_1 _6420_ (.A(_1266_),
    .B(_1330_),
    .X(_1450_));
 sky130_fd_sc_hd__xnor2_1 _6421_ (.A(_1450_),
    .B(_1332_),
    .Y(_1451_));
 sky130_fd_sc_hd__and2_1 _6422_ (.A(_1449_),
    .B(_1451_),
    .X(_1452_));
 sky130_fd_sc_hd__xor2_1 _6423_ (.A(_1364_),
    .B(_1428_),
    .X(_1453_));
 sky130_fd_sc_hd__xnor2_1 _6424_ (.A(_1329_),
    .B(_1269_),
    .Y(_1454_));
 sky130_fd_sc_hd__and2_1 _6425_ (.A(_1453_),
    .B(_1454_),
    .X(_1455_));
 sky130_fd_sc_hd__o21ai_1 _6426_ (.A1(_1363_),
    .A2(_1367_),
    .B1(_1365_),
    .Y(_1456_));
 sky130_fd_sc_hd__nor2_1 _6427_ (.A(_1368_),
    .B(_1426_),
    .Y(_1457_));
 sky130_fd_sc_hd__xnor2_1 _6428_ (.A(_1456_),
    .B(_1457_),
    .Y(_1458_));
 sky130_fd_sc_hd__o21ai_1 _6429_ (.A1(_1267_),
    .A2(_1272_),
    .B1(_1270_),
    .Y(_1459_));
 sky130_fd_sc_hd__nor2_1 _6430_ (.A(_1273_),
    .B(_1327_),
    .Y(_1460_));
 sky130_fd_sc_hd__xnor2_1 _6431_ (.A(_1459_),
    .B(_1460_),
    .Y(_1461_));
 sky130_fd_sc_hd__or2_1 _6432_ (.A(_1458_),
    .B(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__xnor2_1 _6433_ (.A(_1369_),
    .B(_1425_),
    .Y(_1463_));
 sky130_fd_sc_hd__xnor2_1 _6434_ (.A(_1274_),
    .B(_1326_),
    .Y(_1464_));
 sky130_fd_sc_hd__or2_1 _6435_ (.A(_1463_),
    .B(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__o21a_1 _6436_ (.A1(_1366_),
    .A2(_1371_),
    .B1(_1370_),
    .X(_1466_));
 sky130_fd_sc_hd__xnor2_1 _6437_ (.A(_1466_),
    .B(_1424_),
    .Y(_1467_));
 sky130_fd_sc_hd__o21a_1 _6438_ (.A1(_1271_),
    .A2(_1277_),
    .B1(_1275_),
    .X(_1468_));
 sky130_fd_sc_hd__xnor2_1 _6439_ (.A(_1468_),
    .B(_1325_),
    .Y(_1469_));
 sky130_fd_sc_hd__nor2_1 _6440_ (.A(_1467_),
    .B(_1469_),
    .Y(_1470_));
 sky130_fd_sc_hd__xnor2_1 _6441_ (.A(_1374_),
    .B(_1423_),
    .Y(_1471_));
 sky130_fd_sc_hd__xor2_1 _6442_ (.A(_1279_),
    .B(_1323_),
    .X(_1472_));
 sky130_fd_sc_hd__nor2_1 _6443_ (.A(_1471_),
    .B(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__inv_2 _6444_ (.A(_1280_),
    .Y(_1474_));
 sky130_fd_sc_hd__nand2_1 _6445_ (.A(_1322_),
    .B(_1474_),
    .Y(_1475_));
 sky130_fd_sc_hd__xor2_1 _6446_ (.A(_1321_),
    .B(_1475_),
    .X(_1476_));
 sky130_fd_sc_hd__and2b_1 _6447_ (.A_N(_1375_),
    .B(_1422_),
    .X(_1477_));
 sky130_fd_sc_hd__xnor2_1 _6448_ (.A(_1421_),
    .B(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__nor2_1 _6449_ (.A(_1476_),
    .B(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__a21bo_1 _6450_ (.A1(_1349_),
    .A2(_1376_),
    .B1_N(_1377_),
    .X(_1480_));
 sky130_fd_sc_hd__xor2_1 _6451_ (.A(_1480_),
    .B(_1420_),
    .X(_1481_));
 sky130_fd_sc_hd__xor2_1 _6452_ (.A(_1283_),
    .B(_1320_),
    .X(_1482_));
 sky130_fd_sc_hd__or2b_1 _6453_ (.A(_1481_),
    .B_N(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__or2_1 _6454_ (.A(_1319_),
    .B(_1284_),
    .X(_1484_));
 sky130_fd_sc_hd__xnor2_1 _6455_ (.A(_1318_),
    .B(_1484_),
    .Y(_1485_));
 sky130_fd_sc_hd__or2b_1 _6456_ (.A(_1378_),
    .B_N(_1419_),
    .X(_1486_));
 sky130_fd_sc_hd__xnor2_1 _6457_ (.A(_1418_),
    .B(_1486_),
    .Y(_1487_));
 sky130_fd_sc_hd__and2_1 _6458_ (.A(_1485_),
    .B(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__a21bo_1 _6459_ (.A1(_1379_),
    .A2(_1380_),
    .B1_N(_1417_),
    .X(_1489_));
 sky130_fd_sc_hd__xnor2_1 _6460_ (.A(_1416_),
    .B(_1489_),
    .Y(_1490_));
 sky130_fd_sc_hd__a21o_1 _6461_ (.A1(_1285_),
    .A2(_1316_),
    .B1(_1315_),
    .X(_1491_));
 sky130_fd_sc_hd__and3_1 _6462_ (.A(_1317_),
    .B(_1490_),
    .C(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__inv_2 _6463_ (.A(_1415_),
    .Y(_1493_));
 sky130_fd_sc_hd__a211o_1 _6464_ (.A1(_1381_),
    .A2(_1493_),
    .B1(_1414_),
    .C1(_1384_),
    .X(_1494_));
 sky130_fd_sc_hd__o211ai_1 _6465_ (.A1(_1384_),
    .A2(_1414_),
    .B1(_1493_),
    .C1(_1381_),
    .Y(_1495_));
 sky130_fd_sc_hd__nand2_1 _6466_ (.A(_1494_),
    .B(_1495_),
    .Y(_1496_));
 sky130_fd_sc_hd__o21ai_1 _6467_ (.A1(_1313_),
    .A2(_1287_),
    .B1(_1286_),
    .Y(_1497_));
 sky130_fd_sc_hd__nor2_1 _6468_ (.A(_1289_),
    .B(_1312_),
    .Y(_1498_));
 sky130_fd_sc_hd__xnor2_1 _6469_ (.A(_1497_),
    .B(_1498_),
    .Y(_1499_));
 sky130_fd_sc_hd__nor2_1 _6470_ (.A(_1496_),
    .B(_1499_),
    .Y(_1500_));
 sky130_fd_sc_hd__xnor2_1 _6471_ (.A(_1385_),
    .B(_1413_),
    .Y(_1501_));
 sky130_fd_sc_hd__and2_1 _6472_ (.A(_1290_),
    .B(_1311_),
    .X(_1502_));
 sky130_fd_sc_hd__or2_1 _6473_ (.A(_1312_),
    .B(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__nor2_1 _6474_ (.A(_1501_),
    .B(_1503_),
    .Y(_1504_));
 sky130_fd_sc_hd__o21a_1 _6475_ (.A1(_1382_),
    .A2(_1409_),
    .B1(_1386_),
    .X(_1505_));
 sky130_fd_sc_hd__xnor2_1 _6476_ (.A(_1505_),
    .B(_1412_),
    .Y(_1506_));
 sky130_fd_sc_hd__o21a_1 _6477_ (.A1(_1288_),
    .A2(_1307_),
    .B1(_1291_),
    .X(_1507_));
 sky130_fd_sc_hd__xnor2_1 _6478_ (.A(_1507_),
    .B(_1310_),
    .Y(_1508_));
 sky130_fd_sc_hd__nor2_1 _6479_ (.A(_1506_),
    .B(_1508_),
    .Y(_1509_));
 sky130_fd_sc_hd__xor2_1 _6480_ (.A(_1408_),
    .B(_1411_),
    .X(_1510_));
 sky130_fd_sc_hd__xor2_1 _6481_ (.A(_1306_),
    .B(_1309_),
    .X(_1511_));
 sky130_fd_sc_hd__and2_1 _6482_ (.A(_1510_),
    .B(_1511_),
    .X(_1512_));
 sky130_fd_sc_hd__a211oi_1 _6483_ (.A1(_1405_),
    .A2(_1406_),
    .B1(_1389_),
    .C1(_1404_),
    .Y(_1513_));
 sky130_fd_sc_hd__or2_1 _6484_ (.A(_1407_),
    .B(_1513_),
    .X(_1514_));
 sky130_fd_sc_hd__a211oi_1 _6485_ (.A1(_1303_),
    .A2(_1304_),
    .B1(_1294_),
    .C1(_1302_),
    .Y(_1515_));
 sky130_fd_sc_hd__or2_1 _6486_ (.A(_1305_),
    .B(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__nor2_1 _6487_ (.A(_1514_),
    .B(_1516_),
    .Y(_1517_));
 sky130_fd_sc_hd__or3b_1 _6488_ (.A(_1390_),
    .B(_1401_),
    .C_N(_1403_),
    .X(_1518_));
 sky130_fd_sc_hd__nor2b_1 _6489_ (.A(_1404_),
    .B_N(_1518_),
    .Y(_1519_));
 sky130_fd_sc_hd__nor3b_1 _6490_ (.A(_1295_),
    .B(_1299_),
    .C_N(_1301_),
    .Y(_1520_));
 sky130_fd_sc_hd__nor2_1 _6491_ (.A(_1302_),
    .B(_1520_),
    .Y(_1521_));
 sky130_fd_sc_hd__and2_1 _6492_ (.A(_1519_),
    .B(_1521_),
    .X(_1522_));
 sky130_fd_sc_hd__a211o_1 _6493_ (.A1(_1399_),
    .A2(_1400_),
    .B1(_1391_),
    .C1(_1398_),
    .X(_1523_));
 sky130_fd_sc_hd__nand2b_1 _6494_ (.A_N(_1401_),
    .B(_1523_),
    .Y(_1524_));
 sky130_fd_sc_hd__a21oi_1 _6495_ (.A1(_1296_),
    .A2(_1297_),
    .B1(_1298_),
    .Y(_1525_));
 sky130_fd_sc_hd__or2_1 _6496_ (.A(_1299_),
    .B(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__nor2_1 _6497_ (.A(_1524_),
    .B(_1526_),
    .Y(_1527_));
 sky130_fd_sc_hd__nand2_1 _6498_ (.A(_1392_),
    .B(_1393_),
    .Y(_1528_));
 sky130_fd_sc_hd__xor2_1 _6499_ (.A(_1528_),
    .B(_1397_),
    .X(_1529_));
 sky130_fd_sc_hd__nand4_1 _6500_ (.A(_3503_),
    .B(_3536_),
    .C(_1251_),
    .D(_1255_),
    .Y(_1530_));
 sky130_fd_sc_hd__and3_1 _6501_ (.A(_3586_),
    .B(_3503_),
    .C(_1255_),
    .X(_1531_));
 sky130_fd_sc_hd__a22o_1 _6502_ (.A1(_3503_),
    .A2(_1251_),
    .B1(_1255_),
    .B2(_3586_),
    .X(_1532_));
 sky130_fd_sc_hd__a21bo_1 _6503_ (.A1(_1251_),
    .A2(_1531_),
    .B1_N(_1532_),
    .X(_1533_));
 sky130_fd_sc_hd__xnor2_1 _6504_ (.A(_1530_),
    .B(_1533_),
    .Y(_1534_));
 sky130_fd_sc_hd__nor2_1 _6505_ (.A(_1529_),
    .B(_1534_),
    .Y(_1535_));
 sky130_fd_sc_hd__a22o_1 _6506_ (.A1(_3536_),
    .A2(_1251_),
    .B1(_1255_),
    .B2(_3503_),
    .X(_1536_));
 sky130_fd_sc_hd__nor2_1 _6507_ (.A(_1394_),
    .B(_1395_),
    .Y(_1537_));
 sky130_fd_sc_hd__a22oi_1 _6508_ (.A1(_3576_),
    .A2(\M1.U1.U3.u2.instance13_12.Prop_L ),
    .B1(_1352_),
    .B2(_3426_),
    .Y(_1538_));
 sky130_fd_sc_hd__nor2_1 _6509_ (.A(_1396_),
    .B(_1538_),
    .Y(_1539_));
 sky130_fd_sc_hd__xnor2_1 _6510_ (.A(_1537_),
    .B(_1539_),
    .Y(_1540_));
 sky130_fd_sc_hd__and3_1 _6511_ (.A(_1530_),
    .B(_1536_),
    .C(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__a21oi_1 _6512_ (.A1(_1530_),
    .A2(_1536_),
    .B1(_1540_),
    .Y(_1542_));
 sky130_fd_sc_hd__or2_1 _6513_ (.A(_1541_),
    .B(_1542_),
    .X(_1543_));
 sky130_fd_sc_hd__and2_1 _6514_ (.A(_3503_),
    .B(_1347_),
    .X(_1544_));
 sky130_fd_sc_hd__a21o_1 _6515_ (.A1(_3586_),
    .A2(_1352_),
    .B1(_1544_),
    .X(_1545_));
 sky130_fd_sc_hd__and2_1 _6516_ (.A(_3536_),
    .B(_1352_),
    .X(_1546_));
 sky130_fd_sc_hd__and3_1 _6517_ (.A(_1544_),
    .B(_1546_),
    .C(_1395_),
    .X(_1547_));
 sky130_fd_sc_hd__a21o_1 _6518_ (.A1(_1537_),
    .A2(_1545_),
    .B1(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__and3_1 _6519_ (.A(_3546_),
    .B(_1255_),
    .C(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__nor2b_1 _6520_ (.A(_1543_),
    .B_N(_1549_),
    .Y(_1550_));
 sky130_fd_sc_hd__and2_1 _6521_ (.A(_1529_),
    .B(_1534_),
    .X(_1551_));
 sky130_fd_sc_hd__nor2_1 _6522_ (.A(_1535_),
    .B(_1551_),
    .Y(_1552_));
 sky130_fd_sc_hd__o21a_1 _6523_ (.A1(_1541_),
    .A2(_1550_),
    .B1(_1552_),
    .X(_1553_));
 sky130_fd_sc_hd__and2_1 _6524_ (.A(_1524_),
    .B(_1526_),
    .X(_1554_));
 sky130_fd_sc_hd__nor2_1 _6525_ (.A(_1527_),
    .B(_1554_),
    .Y(_1555_));
 sky130_fd_sc_hd__o21a_1 _6526_ (.A1(_1535_),
    .A2(_1553_),
    .B1(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__nor2_1 _6527_ (.A(_1519_),
    .B(_1521_),
    .Y(_1557_));
 sky130_fd_sc_hd__nor2_1 _6528_ (.A(_1522_),
    .B(_1557_),
    .Y(_1558_));
 sky130_fd_sc_hd__o21a_1 _6529_ (.A1(_1527_),
    .A2(_1556_),
    .B1(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__and2_1 _6530_ (.A(_1514_),
    .B(_1516_),
    .X(_1560_));
 sky130_fd_sc_hd__nor2_1 _6531_ (.A(_1517_),
    .B(_1560_),
    .Y(_1561_));
 sky130_fd_sc_hd__o21a_1 _6532_ (.A1(_1522_),
    .A2(_1559_),
    .B1(_1561_),
    .X(_1562_));
 sky130_fd_sc_hd__nor2_1 _6533_ (.A(_1510_),
    .B(_1511_),
    .Y(_1563_));
 sky130_fd_sc_hd__nor2_1 _6534_ (.A(_1512_),
    .B(_1563_),
    .Y(_1564_));
 sky130_fd_sc_hd__o21a_1 _6535_ (.A1(_1517_),
    .A2(_1562_),
    .B1(_1564_),
    .X(_1565_));
 sky130_fd_sc_hd__and2_1 _6536_ (.A(_1506_),
    .B(_1508_),
    .X(_1566_));
 sky130_fd_sc_hd__nor2_1 _6537_ (.A(_1509_),
    .B(_1566_),
    .Y(_1567_));
 sky130_fd_sc_hd__o21a_1 _6538_ (.A1(_1512_),
    .A2(_1565_),
    .B1(_1567_),
    .X(_1568_));
 sky130_fd_sc_hd__and2_1 _6539_ (.A(_1501_),
    .B(_1503_),
    .X(_1569_));
 sky130_fd_sc_hd__nor2_1 _6540_ (.A(_1504_),
    .B(_1569_),
    .Y(_1570_));
 sky130_fd_sc_hd__o21a_1 _6541_ (.A1(_1509_),
    .A2(_1568_),
    .B1(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__xor2_1 _6542_ (.A(_1496_),
    .B(_1499_),
    .X(_1572_));
 sky130_fd_sc_hd__o21a_1 _6543_ (.A1(_1504_),
    .A2(_1571_),
    .B1(_1572_),
    .X(_1573_));
 sky130_fd_sc_hd__a21oi_1 _6544_ (.A1(_1317_),
    .A2(_1491_),
    .B1(_1490_),
    .Y(_1574_));
 sky130_fd_sc_hd__nor2_1 _6545_ (.A(_1492_),
    .B(_1574_),
    .Y(_1575_));
 sky130_fd_sc_hd__o21a_1 _6546_ (.A1(_1500_),
    .A2(_1573_),
    .B1(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__nor2_1 _6547_ (.A(_1485_),
    .B(_1487_),
    .Y(_1577_));
 sky130_fd_sc_hd__or2_1 _6548_ (.A(_1488_),
    .B(_1577_),
    .X(_1578_));
 sky130_fd_sc_hd__o21ba_1 _6549_ (.A1(_1492_),
    .A2(_1576_),
    .B1_N(_1578_),
    .X(_1579_));
 sky130_fd_sc_hd__xnor2_1 _6550_ (.A(_1481_),
    .B(_1482_),
    .Y(_1580_));
 sky130_fd_sc_hd__o21ai_1 _6551_ (.A1(_1488_),
    .A2(_1579_),
    .B1(_1580_),
    .Y(_1581_));
 sky130_fd_sc_hd__nand2_1 _6552_ (.A(_1476_),
    .B(_1478_),
    .Y(_1582_));
 sky130_fd_sc_hd__nand2b_1 _6553_ (.A_N(_1479_),
    .B(_1582_),
    .Y(_1583_));
 sky130_fd_sc_hd__a21oi_1 _6554_ (.A1(_1483_),
    .A2(_1581_),
    .B1(_1583_),
    .Y(_1584_));
 sky130_fd_sc_hd__and2_1 _6555_ (.A(_1471_),
    .B(_1472_),
    .X(_1585_));
 sky130_fd_sc_hd__nor2_1 _6556_ (.A(_1473_),
    .B(_1585_),
    .Y(_1586_));
 sky130_fd_sc_hd__o21a_1 _6557_ (.A1(_1479_),
    .A2(_1584_),
    .B1(_1586_),
    .X(_1587_));
 sky130_fd_sc_hd__and2_1 _6558_ (.A(_1467_),
    .B(_1469_),
    .X(_1588_));
 sky130_fd_sc_hd__nor2_1 _6559_ (.A(_1470_),
    .B(_1588_),
    .Y(_1589_));
 sky130_fd_sc_hd__o21a_1 _6560_ (.A1(_1473_),
    .A2(_1587_),
    .B1(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__nand2_1 _6561_ (.A(_1463_),
    .B(_1464_),
    .Y(_1591_));
 sky130_fd_sc_hd__and2_1 _6562_ (.A(_1465_),
    .B(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__o21ai_1 _6563_ (.A1(_1470_),
    .A2(_1590_),
    .B1(_1592_),
    .Y(_1593_));
 sky130_fd_sc_hd__xnor2_1 _6564_ (.A(_1458_),
    .B(_1461_),
    .Y(_1594_));
 sky130_fd_sc_hd__a21o_1 _6565_ (.A1(_1465_),
    .A2(_1593_),
    .B1(_1594_),
    .X(_1595_));
 sky130_fd_sc_hd__nor2_1 _6566_ (.A(_1453_),
    .B(_1454_),
    .Y(_1596_));
 sky130_fd_sc_hd__or2_1 _6567_ (.A(_1455_),
    .B(_1596_),
    .X(_1597_));
 sky130_fd_sc_hd__a21oi_1 _6568_ (.A1(_1462_),
    .A2(_1595_),
    .B1(_1597_),
    .Y(_1598_));
 sky130_fd_sc_hd__xnor2_1 _6569_ (.A(_1449_),
    .B(_1451_),
    .Y(_1599_));
 sky130_fd_sc_hd__o21ba_1 _6570_ (.A1(_1455_),
    .A2(_1598_),
    .B1_N(_1599_),
    .X(_1600_));
 sky130_fd_sc_hd__xor2_1 _6571_ (.A(_1444_),
    .B(_1446_),
    .X(_1601_));
 sky130_fd_sc_hd__o21a_1 _6572_ (.A1(_1452_),
    .A2(_1600_),
    .B1(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__xor2_1 _6573_ (.A(_1440_),
    .B(_1441_),
    .X(_1603_));
 sky130_fd_sc_hd__o21a_1 _6574_ (.A1(_1447_),
    .A2(_1602_),
    .B1(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__xnor2_1 _6575_ (.A(_1435_),
    .B(_1437_),
    .Y(_1605_));
 sky130_fd_sc_hd__o21ba_1 _6576_ (.A1(_1442_),
    .A2(_1604_),
    .B1_N(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__nand2_1 _6577_ (.A(_1350_),
    .B(_1434_),
    .Y(_1607_));
 sky130_fd_sc_hd__xor2_1 _6578_ (.A(_1351_),
    .B(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__o21ba_1 _6579_ (.A1(_1438_),
    .A2(_1606_),
    .B1_N(_1608_),
    .X(_1609_));
 sky130_fd_sc_hd__a31o_1 _6580_ (.A1(_1350_),
    .A2(_1351_),
    .A3(_1434_),
    .B1(_1609_),
    .X(_1610_));
 sky130_fd_sc_hd__nand2_1 _6581_ (.A(_1346_),
    .B(_1610_),
    .Y(_1611_));
 sky130_fd_sc_hd__nor2_1 _6582_ (.A(_1438_),
    .B(_1606_),
    .Y(_1612_));
 sky130_fd_sc_hd__xnor2_1 _6583_ (.A(_1608_),
    .B(_1612_),
    .Y(_1613_));
 sky130_fd_sc_hd__nor2_1 _6584_ (.A(_1442_),
    .B(_1604_),
    .Y(_1614_));
 sky130_fd_sc_hd__and2_1 _6585_ (.A(_1605_),
    .B(_1614_),
    .X(_1615_));
 sky130_fd_sc_hd__or2_1 _6586_ (.A(_1606_),
    .B(_1615_),
    .X(_1616_));
 sky130_fd_sc_hd__buf_2 _6587_ (.A(\M1.U1.U2.u2.instance11_10.Prop_L ),
    .X(_1617_));
 sky130_fd_sc_hd__clkbuf_2 _6588_ (.A(_1617_),
    .X(_1618_));
 sky130_fd_sc_hd__clkbuf_2 _6589_ (.A(_1618_),
    .X(_1619_));
 sky130_fd_sc_hd__buf_2 _6590_ (.A(_1619_),
    .X(_1620_));
 sky130_fd_sc_hd__buf_6 _6591_ (.A(\M1.U1.U1.u2.instance9_8.Prop_L ),
    .X(_1621_));
 sky130_fd_sc_hd__buf_6 _6592_ (.A(_1621_),
    .X(_1622_));
 sky130_fd_sc_hd__clkbuf_2 _6593_ (.A(_1622_),
    .X(_1623_));
 sky130_fd_sc_hd__buf_2 _6594_ (.A(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__clkbuf_2 _6595_ (.A(_1624_),
    .X(_1625_));
 sky130_fd_sc_hd__buf_6 _6596_ (.A(\In2_reg[0] ),
    .X(_1626_));
 sky130_fd_sc_hd__buf_2 _6597_ (.A(_1626_),
    .X(_1627_));
 sky130_fd_sc_hd__clkbuf_2 _6598_ (.A(_1627_),
    .X(_1628_));
 sky130_fd_sc_hd__buf_2 _6599_ (.A(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__and4_1 _6600_ (.A(\In1_reg[21] ),
    .B(_2557_),
    .C(_1625_),
    .D(_1629_),
    .X(_1630_));
 sky130_fd_sc_hd__and4_1 _6601_ (.A(\In1_reg[20] ),
    .B(_2612_),
    .C(_1625_),
    .D(_1629_),
    .X(_1631_));
 sky130_fd_sc_hd__nand2_1 _6602_ (.A(\In1_reg[19] ),
    .B(_1624_),
    .Y(_1632_));
 sky130_fd_sc_hd__nand2_1 _6603_ (.A(\In1_reg[18] ),
    .B(_1628_),
    .Y(_1633_));
 sky130_fd_sc_hd__nor2_1 _6604_ (.A(_1632_),
    .B(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__nand2_1 _6605_ (.A(\In1_reg[17] ),
    .B(_1624_),
    .Y(_1635_));
 sky130_fd_sc_hd__and4_1 _6606_ (.A(\In1_reg[18] ),
    .B(\In1_reg[17] ),
    .C(_1624_),
    .D(_1628_),
    .X(_1636_));
 sky130_fd_sc_hd__a21o_1 _6607_ (.A1(_1633_),
    .A2(_1635_),
    .B1(_1636_),
    .X(_1637_));
 sky130_fd_sc_hd__inv_2 _6608_ (.A(_1637_),
    .Y(_1638_));
 sky130_fd_sc_hd__nand2_1 _6609_ (.A(\In1_reg[16] ),
    .B(_1628_),
    .Y(_1639_));
 sky130_fd_sc_hd__nor2_1 _6610_ (.A(_1635_),
    .B(_1639_),
    .Y(_1640_));
 sky130_fd_sc_hd__a22o_1 _6611_ (.A1(_2854_),
    .A2(_1624_),
    .B1(_1628_),
    .B2(\In1_reg[15] ),
    .X(_1641_));
 sky130_fd_sc_hd__and4_1 _6612_ (.A(\In1_reg[13] ),
    .B(\In1_reg[12] ),
    .C(_1623_),
    .D(_1628_),
    .X(_1642_));
 sky130_fd_sc_hd__and4_1 _6613_ (.A(\In1_reg[12] ),
    .B(_3019_),
    .C(_1623_),
    .D(_1627_),
    .X(_1643_));
 sky130_fd_sc_hd__and4_1 _6614_ (.A(\In1_reg[11] ),
    .B(\In1_reg[10] ),
    .C(_1623_),
    .D(_1627_),
    .X(_1644_));
 sky130_fd_sc_hd__and4_1 _6615_ (.A(_3074_),
    .B(_3118_),
    .C(_1623_),
    .D(_1627_),
    .X(_1645_));
 sky130_fd_sc_hd__and4_1 _6616_ (.A(\In1_reg[9] ),
    .B(\In1_reg[8] ),
    .C(_1622_),
    .D(_1626_),
    .X(_1646_));
 sky130_fd_sc_hd__and4_1 _6617_ (.A(\In1_reg[8] ),
    .B(\In1_reg[7] ),
    .C(_1622_),
    .D(_1626_),
    .X(_1647_));
 sky130_fd_sc_hd__and4_1 _6618_ (.A(\In1_reg[6] ),
    .B(\In1_reg[5] ),
    .C(_1621_),
    .D(\In2_reg[0] ),
    .X(_1648_));
 sky130_fd_sc_hd__and4_1 _6619_ (.A(\In1_reg[7] ),
    .B(\In1_reg[6] ),
    .C(_1621_),
    .D(\In2_reg[0] ),
    .X(_1649_));
 sky130_fd_sc_hd__and3_1 _6620_ (.A(\In1_reg[5] ),
    .B(\In1_reg[4] ),
    .C(\In2_reg[0] ),
    .X(_1650_));
 sky130_fd_sc_hd__and4_1 _6621_ (.A(\In2_reg[0] ),
    .B(\In1_reg[3] ),
    .C(\M1.U1.U1.u2.instance9_8.Prop_L ),
    .D(\In1_reg[4] ),
    .X(_1651_));
 sky130_fd_sc_hd__a21oi_1 _6622_ (.A1(_1622_),
    .A2(_1650_),
    .B1(_1651_),
    .Y(_1652_));
 sky130_fd_sc_hd__a22o_1 _6623_ (.A1(\In1_reg[3] ),
    .A2(_1621_),
    .B1(\In2_reg[0] ),
    .B2(\In1_reg[4] ),
    .X(_1653_));
 sky130_fd_sc_hd__nand2b_2 _6624_ (.A_N(_1651_),
    .B(_1653_),
    .Y(_1654_));
 sky130_fd_sc_hd__a22o_1 _6625_ (.A1(\In1_reg[4] ),
    .A2(_1621_),
    .B1(\In2_reg[0] ),
    .B2(\In1_reg[5] ),
    .X(_1655_));
 sky130_fd_sc_hd__and4_1 _6626_ (.A(net126),
    .B(_3536_),
    .C(_1621_),
    .D(\In2_reg[0] ),
    .X(_1656_));
 sky130_fd_sc_hd__o2111a_1 _6627_ (.A1(\In1_reg[3] ),
    .A2(\In1_reg[1] ),
    .B1(_1621_),
    .C1(\In2_reg[0] ),
    .D1(_3576_),
    .X(_1657_));
 sky130_fd_sc_hd__a21o_4 _6628_ (.A1(_1656_),
    .A2(_3426_),
    .B1(_1657_),
    .X(_1658_));
 sky130_fd_sc_hd__nand3b_4 _6629_ (.A_N(_1654_),
    .B(_1655_),
    .C(_1658_),
    .Y(_1659_));
 sky130_fd_sc_hd__a22oi_1 _6630_ (.A1(\In1_reg[5] ),
    .A2(_1621_),
    .B1(_1626_),
    .B2(_3283_),
    .Y(_1660_));
 sky130_fd_sc_hd__or2_1 _6631_ (.A(_1648_),
    .B(_1660_),
    .X(_1661_));
 sky130_fd_sc_hd__a22oi_1 _6632_ (.A1(_3283_),
    .A2(_1621_),
    .B1(_1626_),
    .B2(\In1_reg[7] ),
    .Y(_1662_));
 sky130_fd_sc_hd__or2_1 _6633_ (.A(_1649_),
    .B(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__a211oi_2 _6634_ (.A1(_1652_),
    .A2(_1659_),
    .B1(_1661_),
    .C1(_1663_),
    .Y(_1664_));
 sky130_fd_sc_hd__a22o_1 _6635_ (.A1(\In1_reg[7] ),
    .A2(_1622_),
    .B1(_1627_),
    .B2(\In1_reg[8] ),
    .X(_1665_));
 sky130_fd_sc_hd__inv_2 _6636_ (.A(_1647_),
    .Y(_1666_));
 sky130_fd_sc_hd__o311a_1 _6637_ (.A1(_1648_),
    .A2(_1664_),
    .A3(_1649_),
    .B1(_1665_),
    .C1(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__inv_4 _6638_ (.A(_1646_),
    .Y(_1668_));
 sky130_fd_sc_hd__a22o_1 _6639_ (.A1(\In1_reg[8] ),
    .A2(_1622_),
    .B1(_1627_),
    .B2(\In1_reg[9] ),
    .X(_1669_));
 sky130_fd_sc_hd__o211a_1 _6640_ (.A1(_1667_),
    .A2(_1647_),
    .B1(_1668_),
    .C1(_1669_),
    .X(_1670_));
 sky130_fd_sc_hd__a22o_1 _6641_ (.A1(\In1_reg[9] ),
    .A2(_1623_),
    .B1(_1627_),
    .B2(\In1_reg[10] ),
    .X(_1671_));
 sky130_fd_sc_hd__nand4_1 _6642_ (.A(\In1_reg[10] ),
    .B(_3118_),
    .C(_1623_),
    .D(_1627_),
    .Y(_1672_));
 sky130_fd_sc_hd__o211a_1 _6643_ (.A1(_1670_),
    .A2(_1646_),
    .B1(_1671_),
    .C1(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__a22oi_1 _6644_ (.A1(\In1_reg[10] ),
    .A2(_1623_),
    .B1(_1627_),
    .B2(\In1_reg[11] ),
    .Y(_1674_));
 sky130_fd_sc_hd__nor2_1 _6645_ (.A(_1644_),
    .B(_1674_),
    .Y(_1675_));
 sky130_fd_sc_hd__o21a_1 _6646_ (.A1(_1673_),
    .A2(_1645_),
    .B1(_1675_),
    .X(_1677_));
 sky130_fd_sc_hd__a22oi_1 _6647_ (.A1(_3019_),
    .A2(_1623_),
    .B1(_1627_),
    .B2(\In1_reg[12] ),
    .Y(_1678_));
 sky130_fd_sc_hd__nor2_1 _6648_ (.A(_1643_),
    .B(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__o21a_1 _6649_ (.A1(_1677_),
    .A2(_1644_),
    .B1(_1679_),
    .X(_1680_));
 sky130_fd_sc_hd__a22oi_1 _6650_ (.A1(\In1_reg[12] ),
    .A2(_1624_),
    .B1(_1628_),
    .B2(\In1_reg[13] ),
    .Y(_1681_));
 sky130_fd_sc_hd__nor2_1 _6651_ (.A(_1642_),
    .B(_1681_),
    .Y(_1682_));
 sky130_fd_sc_hd__o21a_1 _6652_ (.A1(_1680_),
    .A2(_1643_),
    .B1(_1682_),
    .X(_1683_));
 sky130_fd_sc_hd__nand2_1 _6653_ (.A(_2898_),
    .B(_1624_),
    .Y(_1684_));
 sky130_fd_sc_hd__nand2_1 _6654_ (.A(\In1_reg[14] ),
    .B(_1628_),
    .Y(_1685_));
 sky130_fd_sc_hd__and4_1 _6655_ (.A(\In1_reg[14] ),
    .B(\In1_reg[13] ),
    .C(_1623_),
    .D(_1628_),
    .X(_1686_));
 sky130_fd_sc_hd__a21o_1 _6656_ (.A1(_1684_),
    .A2(_1685_),
    .B1(_1686_),
    .X(_1688_));
 sky130_fd_sc_hd__o21ba_4 _6657_ (.A1(_1642_),
    .A2(_1683_),
    .B1_N(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__nand2_1 _6658_ (.A(\In1_reg[15] ),
    .B(_1624_),
    .Y(_1690_));
 sky130_fd_sc_hd__nor2_1 _6659_ (.A(_1685_),
    .B(_1690_),
    .Y(_1691_));
 sky130_fd_sc_hd__a211o_1 _6660_ (.A1(_1689_),
    .A2(_1641_),
    .B1(_1691_),
    .C1(_1686_),
    .X(_1692_));
 sky130_fd_sc_hd__and4_1 _6661_ (.A(\In1_reg[16] ),
    .B(\In1_reg[15] ),
    .C(_1624_),
    .D(_1628_),
    .X(_1693_));
 sky130_fd_sc_hd__a21oi_1 _6662_ (.A1(_1639_),
    .A2(_1690_),
    .B1(_1693_),
    .Y(_1694_));
 sky130_fd_sc_hd__a21o_1 _6663_ (.A1(_1694_),
    .A2(_1692_),
    .B1(_1693_),
    .X(_1695_));
 sky130_fd_sc_hd__a22o_1 _6664_ (.A1(\In1_reg[16] ),
    .A2(_1624_),
    .B1(_1629_),
    .B2(\In1_reg[17] ),
    .X(_1696_));
 sky130_fd_sc_hd__o21a_1 _6665_ (.A1(_1695_),
    .A2(_1640_),
    .B1(_1696_),
    .X(_1697_));
 sky130_fd_sc_hd__a21o_1 _6666_ (.A1(_1697_),
    .A2(_1638_),
    .B1(_1636_),
    .X(_1698_));
 sky130_fd_sc_hd__a21boi_1 _6667_ (.A1(_2557_),
    .A2(_1629_),
    .B1_N(_1632_),
    .Y(_1699_));
 sky130_fd_sc_hd__nor2_1 _6668_ (.A(_1631_),
    .B(_1699_),
    .Y(_1700_));
 sky130_fd_sc_hd__a22o_1 _6669_ (.A1(_2667_),
    .A2(_1625_),
    .B1(_1629_),
    .B2(_2612_),
    .X(_1701_));
 sky130_fd_sc_hd__o211a_1 _6670_ (.A1(_1698_),
    .A2(_1634_),
    .B1(_1700_),
    .C1(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__a22oi_1 _6671_ (.A1(_2557_),
    .A2(_1625_),
    .B1(_1629_),
    .B2(_2469_),
    .Y(_1703_));
 sky130_fd_sc_hd__nor2_1 _6672_ (.A(_1630_),
    .B(_1703_),
    .Y(_1704_));
 sky130_fd_sc_hd__o21a_1 _6673_ (.A1(_1702_),
    .A2(_1631_),
    .B1(_1704_),
    .X(_1705_));
 sky130_fd_sc_hd__a22o_1 _6674_ (.A1(_2469_),
    .A2(_1625_),
    .B1(_1629_),
    .B2(\In1_reg[22] ),
    .X(_1706_));
 sky130_fd_sc_hd__nand4_1 _6675_ (.A(\In1_reg[22] ),
    .B(_2469_),
    .C(_1625_),
    .D(_1629_),
    .Y(_1707_));
 sky130_fd_sc_hd__o211a_4 _6676_ (.A1(_1630_),
    .A2(_1705_),
    .B1(_1706_),
    .C1(_1707_),
    .X(_1709_));
 sky130_fd_sc_hd__and3_1 _6677_ (.A(\In1_reg[22] ),
    .B(_1625_),
    .C(_1629_),
    .X(_1710_));
 sky130_fd_sc_hd__or2_1 _6678_ (.A(_1709_),
    .B(_1710_),
    .X(_1711_));
 sky130_fd_sc_hd__buf_2 _6679_ (.A(\In2_reg[2] ),
    .X(_1712_));
 sky130_fd_sc_hd__clkbuf_2 _6680_ (.A(_1712_),
    .X(_1713_));
 sky130_fd_sc_hd__clkbuf_2 _6681_ (.A(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__buf_2 _6682_ (.A(_1714_),
    .X(_1715_));
 sky130_fd_sc_hd__and3_1 _6683_ (.A(_3800_),
    .B(_1620_),
    .C(_1715_),
    .X(_1716_));
 sky130_fd_sc_hd__a21oi_1 _6684_ (.A1(_3800_),
    .A2(_1620_),
    .B1(_1715_),
    .Y(_1717_));
 sky130_fd_sc_hd__or2_1 _6685_ (.A(_1716_),
    .B(_1717_),
    .X(_1718_));
 sky130_fd_sc_hd__a21bo_1 _6686_ (.A1(_2480_),
    .A2(_1715_),
    .B1_N(_1718_),
    .X(_1719_));
 sky130_fd_sc_hd__a22o_1 _6687_ (.A1(_2557_),
    .A2(_1620_),
    .B1(_1715_),
    .B2(_2469_),
    .X(_1720_));
 sky130_fd_sc_hd__nand2_1 _6688_ (.A(_2612_),
    .B(_1620_),
    .Y(_1721_));
 sky130_fd_sc_hd__nand2_1 _6689_ (.A(_2557_),
    .B(_1715_),
    .Y(_1722_));
 sky130_fd_sc_hd__and4_1 _6690_ (.A(_2557_),
    .B(_2612_),
    .C(_1620_),
    .D(_1715_),
    .X(_1723_));
 sky130_fd_sc_hd__a21o_1 _6691_ (.A1(_1721_),
    .A2(_1722_),
    .B1(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__a22o_1 _6692_ (.A1(_2667_),
    .A2(_1620_),
    .B1(_1715_),
    .B2(_2612_),
    .X(_1725_));
 sky130_fd_sc_hd__and4_1 _6693_ (.A(\In1_reg[18] ),
    .B(\In1_reg[17] ),
    .C(_1619_),
    .D(_1714_),
    .X(_1726_));
 sky130_fd_sc_hd__and4_1 _6694_ (.A(_2711_),
    .B(_2777_),
    .C(_1619_),
    .D(_1714_),
    .X(_1727_));
 sky130_fd_sc_hd__and3_1 _6695_ (.A(\In1_reg[16] ),
    .B(\In1_reg[15] ),
    .C(_1714_),
    .X(_1728_));
 sky130_fd_sc_hd__a22o_1 _6696_ (.A1(_2821_),
    .A2(_1619_),
    .B1(_1714_),
    .B2(\In1_reg[16] ),
    .X(_1730_));
 sky130_fd_sc_hd__a21bo_1 _6697_ (.A1(_1619_),
    .A2(_1728_),
    .B1_N(_1730_),
    .X(_1731_));
 sky130_fd_sc_hd__and4_1 _6698_ (.A(_2821_),
    .B(_2854_),
    .C(_1619_),
    .D(_1714_),
    .X(_1732_));
 sky130_fd_sc_hd__and2_1 _6699_ (.A(_2854_),
    .B(_1619_),
    .X(_1733_));
 sky130_fd_sc_hd__and2_1 _6700_ (.A(\In1_reg[13] ),
    .B(_1714_),
    .X(_1734_));
 sky130_fd_sc_hd__a21o_1 _6701_ (.A1(_2975_),
    .A2(_1618_),
    .B1(_1734_),
    .X(_1735_));
 sky130_fd_sc_hd__nand2_1 _6702_ (.A(_3019_),
    .B(_1618_),
    .Y(_1736_));
 sky130_fd_sc_hd__nand2_1 _6703_ (.A(_3074_),
    .B(_1713_),
    .Y(_1737_));
 sky130_fd_sc_hd__or2_1 _6704_ (.A(_1736_),
    .B(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__and4_1 _6705_ (.A(\In1_reg[10] ),
    .B(_3118_),
    .C(_1618_),
    .D(_1713_),
    .X(_1739_));
 sky130_fd_sc_hd__and4_1 _6706_ (.A(\In1_reg[9] ),
    .B(_3162_),
    .C(_1617_),
    .D(_1713_),
    .X(_1740_));
 sky130_fd_sc_hd__and4_1 _6707_ (.A(_3162_),
    .B(_3217_),
    .C(_1618_),
    .D(_1713_),
    .X(_1741_));
 sky130_fd_sc_hd__and4_1 _6708_ (.A(\In1_reg[7] ),
    .B(_3283_),
    .C(_1617_),
    .D(_1712_),
    .X(_1742_));
 sky130_fd_sc_hd__and4_1 _6709_ (.A(\In1_reg[6] ),
    .B(\In1_reg[5] ),
    .C(\M1.U1.U2.u2.instance11_10.Prop_L ),
    .D(_1712_),
    .X(_1743_));
 sky130_fd_sc_hd__and4_1 _6710_ (.A(\M1.U1.U2.u2.instance11_10.Prop_L ),
    .B(\In1_reg[0] ),
    .C(\In1_reg[1] ),
    .D(\In2_reg[2] ),
    .X(_1744_));
 sky130_fd_sc_hd__and4_1 _6711_ (.A(\M1.U1.U2.u2.instance11_10.Prop_L ),
    .B(\In1_reg[2] ),
    .C(\In1_reg[3] ),
    .D(\In2_reg[2] ),
    .X(_1745_));
 sky130_fd_sc_hd__and4_1 _6712_ (.A(\In1_reg[2] ),
    .B(\In1_reg[1] ),
    .C(\M1.U1.U2.u2.instance11_10.Prop_L ),
    .D(\In2_reg[2] ),
    .X(_1746_));
 sky130_fd_sc_hd__a211o_1 _6713_ (.A1(\In1_reg[5] ),
    .A2(_1744_),
    .B1(_1745_),
    .C1(_1746_),
    .X(_1747_));
 sky130_fd_sc_hd__and4_1 _6714_ (.A(\In1_reg[4] ),
    .B(\In1_reg[3] ),
    .C(\M1.U1.U2.u2.instance11_10.Prop_L ),
    .D(\In2_reg[2] ),
    .X(_1748_));
 sky130_fd_sc_hd__a22oi_1 _6715_ (.A1(_3426_),
    .A2(\M1.U1.U2.u2.instance11_10.Prop_L ),
    .B1(\In2_reg[2] ),
    .B2(\In1_reg[4] ),
    .Y(_1749_));
 sky130_fd_sc_hd__nor2_1 _6716_ (.A(_1748_),
    .B(_1749_),
    .Y(_1751_));
 sky130_fd_sc_hd__a22o_1 _6717_ (.A1(\In1_reg[4] ),
    .A2(\M1.U1.U2.u2.instance11_10.Prop_L ),
    .B1(\In2_reg[2] ),
    .B2(\In1_reg[5] ),
    .X(_1752_));
 sky130_fd_sc_hd__and3_1 _6718_ (.A(_1747_),
    .B(_1751_),
    .C(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__nand4_1 _6719_ (.A(_3338_),
    .B(_3380_),
    .C(_1617_),
    .D(_1712_),
    .Y(_1754_));
 sky130_fd_sc_hd__or2b_1 _6720_ (.A(_1748_),
    .B_N(_1754_),
    .X(_1755_));
 sky130_fd_sc_hd__a22o_1 _6721_ (.A1(_3338_),
    .A2(_1617_),
    .B1(_1712_),
    .B2(_3283_),
    .X(_1756_));
 sky130_fd_sc_hd__inv_2 _6722_ (.A(_1743_),
    .Y(_1757_));
 sky130_fd_sc_hd__o211a_1 _6723_ (.A1(_1755_),
    .A2(_1753_),
    .B1(_1756_),
    .C1(_1757_),
    .X(_1758_));
 sky130_fd_sc_hd__inv_2 _6724_ (.A(_1742_),
    .Y(_1759_));
 sky130_fd_sc_hd__a22o_1 _6725_ (.A1(_3283_),
    .A2(_1617_),
    .B1(_1712_),
    .B2(_3217_),
    .X(_1760_));
 sky130_fd_sc_hd__o211a_1 _6726_ (.A1(_1758_),
    .A2(_1743_),
    .B1(_1759_),
    .C1(_1760_),
    .X(_1761_));
 sky130_fd_sc_hd__a22o_1 _6727_ (.A1(_3217_),
    .A2(_1617_),
    .B1(_1713_),
    .B2(_3162_),
    .X(_1762_));
 sky130_fd_sc_hd__nand4_1 _6728_ (.A(_3162_),
    .B(_3217_),
    .C(_1617_),
    .D(_1713_),
    .Y(_1763_));
 sky130_fd_sc_hd__o211a_1 _6729_ (.A1(_1761_),
    .A2(_1742_),
    .B1(_1762_),
    .C1(_1763_),
    .X(_1764_));
 sky130_fd_sc_hd__a22oi_1 _6730_ (.A1(_3162_),
    .A2(_1618_),
    .B1(_1713_),
    .B2(\In1_reg[9] ),
    .Y(_1765_));
 sky130_fd_sc_hd__nor2_1 _6731_ (.A(_1740_),
    .B(_1765_),
    .Y(_1766_));
 sky130_fd_sc_hd__o21a_1 _6732_ (.A1(_1764_),
    .A2(_1741_),
    .B1(_1766_),
    .X(_1767_));
 sky130_fd_sc_hd__nand2_1 _6733_ (.A(_3118_),
    .B(_1618_),
    .Y(_1768_));
 sky130_fd_sc_hd__a21oi_1 _6734_ (.A1(_1737_),
    .A2(_1768_),
    .B1(_1739_),
    .Y(_1769_));
 sky130_fd_sc_hd__o21a_1 _6735_ (.A1(_1767_),
    .A2(_1740_),
    .B1(_1769_),
    .X(_1770_));
 sky130_fd_sc_hd__a22o_1 _6736_ (.A1(_3074_),
    .A2(_1618_),
    .B1(_1713_),
    .B2(_3019_),
    .X(_1772_));
 sky130_fd_sc_hd__o211ai_2 _6737_ (.A1(_1770_),
    .A2(_1739_),
    .B1(_1738_),
    .C1(_1772_),
    .Y(_1773_));
 sky130_fd_sc_hd__nand2_1 _6738_ (.A(_2975_),
    .B(_1714_),
    .Y(_1774_));
 sky130_fd_sc_hd__and4_1 _6739_ (.A(\In1_reg[12] ),
    .B(_3019_),
    .C(_1618_),
    .D(_1713_),
    .X(_1775_));
 sky130_fd_sc_hd__a21o_1 _6740_ (.A1(_1736_),
    .A2(_1774_),
    .B1(_1775_),
    .X(_1776_));
 sky130_fd_sc_hd__a21oi_2 _6741_ (.A1(_1773_),
    .A2(_1738_),
    .B1(_1776_),
    .Y(_1777_));
 sky130_fd_sc_hd__and3_1 _6742_ (.A(_2975_),
    .B(_1618_),
    .C(_1734_),
    .X(_1778_));
 sky130_fd_sc_hd__a211o_1 _6743_ (.A1(_1777_),
    .A2(_1735_),
    .B1(_1778_),
    .C1(_1775_),
    .X(_1779_));
 sky130_fd_sc_hd__a22o_1 _6744_ (.A1(_2898_),
    .A2(_1619_),
    .B1(_1714_),
    .B2(_2854_),
    .X(_1780_));
 sky130_fd_sc_hd__a22o_1 _6745_ (.A1(_1733_),
    .A2(_1734_),
    .B1(_1780_),
    .B2(_1779_),
    .X(_1781_));
 sky130_fd_sc_hd__a21o_1 _6746_ (.A1(_2821_),
    .A2(_1714_),
    .B1(_1733_),
    .X(_1782_));
 sky130_fd_sc_hd__o21ai_2 _6747_ (.A1(_1781_),
    .A2(_1732_),
    .B1(_1782_),
    .Y(_1783_));
 sky130_fd_sc_hd__a2bb2o_4 _6748_ (.A1_N(_1731_),
    .A2_N(_1783_),
    .B1(_1619_),
    .B2(_1728_),
    .X(_1784_));
 sky130_fd_sc_hd__a22o_1 _6749_ (.A1(_2777_),
    .A2(_1620_),
    .B1(_1715_),
    .B2(_2711_),
    .X(_1785_));
 sky130_fd_sc_hd__nand2_1 _6750_ (.A(\In1_reg[18] ),
    .B(_1715_),
    .Y(_1786_));
 sky130_fd_sc_hd__nand2_1 _6751_ (.A(_2711_),
    .B(_1619_),
    .Y(_1787_));
 sky130_fd_sc_hd__a21oi_1 _6752_ (.A1(_1786_),
    .A2(_1787_),
    .B1(_1726_),
    .Y(_1788_));
 sky130_fd_sc_hd__o211a_1 _6753_ (.A1(_1727_),
    .A2(_1784_),
    .B1(_1785_),
    .C1(_1788_),
    .X(_1789_));
 sky130_fd_sc_hd__or2_4 _6754_ (.A(_1726_),
    .B(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__o2bb2a_4 _6755_ (.A1_N(_1725_),
    .A2_N(_1790_),
    .B1(_1721_),
    .B2(_1786_),
    .X(_1791_));
 sky130_fd_sc_hd__nor2_1 _6756_ (.A(_1724_),
    .B(_1791_),
    .Y(_1793_));
 sky130_fd_sc_hd__nand2_1 _6757_ (.A(_2469_),
    .B(_1620_),
    .Y(_1794_));
 sky130_fd_sc_hd__nor2_1 _6758_ (.A(_1722_),
    .B(_1794_),
    .Y(_1795_));
 sky130_fd_sc_hd__a211o_1 _6759_ (.A1(_1793_),
    .A2(_1720_),
    .B1(_1795_),
    .C1(_1723_),
    .X(_1796_));
 sky130_fd_sc_hd__nand2_1 _6760_ (.A(\In1_reg[22] ),
    .B(_1715_),
    .Y(_1797_));
 sky130_fd_sc_hd__xor2_1 _6761_ (.A(_1794_),
    .B(_1797_),
    .X(_1798_));
 sky130_fd_sc_hd__and2_1 _6762_ (.A(_1796_),
    .B(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__mux2_2 _6763_ (.A0(_1719_),
    .A1(_1718_),
    .S(_1799_),
    .X(_1800_));
 sky130_fd_sc_hd__nor2_1 _6764_ (.A(_1709_),
    .B(_1710_),
    .Y(_1801_));
 sky130_fd_sc_hd__xor2_1 _6765_ (.A(_1796_),
    .B(_1798_),
    .X(_1802_));
 sky130_fd_sc_hd__and3_1 _6766_ (.A(_1802_),
    .B(_1801_),
    .C(_1625_),
    .X(_1803_));
 sky130_fd_sc_hd__o21ai_1 _6767_ (.A1(_1722_),
    .A2(_1794_),
    .B1(_1720_),
    .Y(_1804_));
 sky130_fd_sc_hd__nor2_1 _6768_ (.A(_1723_),
    .B(_1793_),
    .Y(_1805_));
 sky130_fd_sc_hd__xnor2_1 _6769_ (.A(_1804_),
    .B(_1805_),
    .Y(_1806_));
 sky130_fd_sc_hd__a21oi_1 _6770_ (.A1(\In1_reg[22] ),
    .A2(_1625_),
    .B1(_1629_),
    .Y(_1807_));
 sky130_fd_sc_hd__or2_1 _6771_ (.A(_1710_),
    .B(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__nand2_1 _6772_ (.A(_1707_),
    .B(_1808_),
    .Y(_1809_));
 sky130_fd_sc_hd__mux2_2 _6773_ (.A0(_1809_),
    .A1(_1808_),
    .S(_1709_),
    .X(_1810_));
 sky130_fd_sc_hd__or2b_1 _6774_ (.A(_1806_),
    .B_N(_1810_),
    .X(_1811_));
 sky130_fd_sc_hd__and2_1 _6775_ (.A(_1724_),
    .B(_1791_),
    .X(_1812_));
 sky130_fd_sc_hd__or2_4 _6776_ (.A(_1793_),
    .B(_1812_),
    .X(_1814_));
 sky130_fd_sc_hd__a211o_1 _6777_ (.A1(_1706_),
    .A2(_1707_),
    .B1(_1705_),
    .C1(_1630_),
    .X(_1815_));
 sky130_fd_sc_hd__or3b_4 _6778_ (.A(_1709_),
    .B(_1814_),
    .C_N(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__nor3_1 _6779_ (.A(_1704_),
    .B(_1631_),
    .C(_1702_),
    .Y(_1817_));
 sky130_fd_sc_hd__o21a_1 _6780_ (.A1(_1721_),
    .A2(_1786_),
    .B1(_1725_),
    .X(_1818_));
 sky130_fd_sc_hd__xnor2_1 _6781_ (.A(_1818_),
    .B(_1790_),
    .Y(_1819_));
 sky130_fd_sc_hd__or3_1 _6782_ (.A(_1705_),
    .B(_1817_),
    .C(_1819_),
    .X(_1820_));
 sky130_fd_sc_hd__o21a_1 _6783_ (.A1(_1634_),
    .A2(_1698_),
    .B1(_1701_),
    .X(_1821_));
 sky130_fd_sc_hd__xnor2_1 _6784_ (.A(_1700_),
    .B(_1821_),
    .Y(_1822_));
 sky130_fd_sc_hd__o21a_1 _6785_ (.A1(_1727_),
    .A2(_1784_),
    .B1(_1785_),
    .X(_1823_));
 sky130_fd_sc_hd__nor2_1 _6786_ (.A(_1788_),
    .B(_1823_),
    .Y(_1824_));
 sky130_fd_sc_hd__or2_1 _6787_ (.A(_1789_),
    .B(_1824_),
    .X(_1825_));
 sky130_fd_sc_hd__nor2_1 _6788_ (.A(_1822_),
    .B(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__and2b_1 _6789_ (.A_N(_1727_),
    .B(_1785_),
    .X(_1827_));
 sky130_fd_sc_hd__xnor2_1 _6790_ (.A(_1784_),
    .B(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__o21a_1 _6791_ (.A1(_1632_),
    .A2(_1633_),
    .B1(_1701_),
    .X(_1829_));
 sky130_fd_sc_hd__xor2_1 _6792_ (.A(_1698_),
    .B(_1829_),
    .X(_1830_));
 sky130_fd_sc_hd__and2b_1 _6793_ (.A_N(_1828_),
    .B(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__xnor2_1 _6794_ (.A(_1637_),
    .B(_1697_),
    .Y(_1832_));
 sky130_fd_sc_hd__xnor2_1 _6795_ (.A(_1731_),
    .B(_1783_),
    .Y(_1833_));
 sky130_fd_sc_hd__inv_2 _6796_ (.A(_1833_),
    .Y(_1835_));
 sky130_fd_sc_hd__or2b_1 _6797_ (.A(_1732_),
    .B_N(_1782_),
    .X(_1836_));
 sky130_fd_sc_hd__xnor2_1 _6798_ (.A(_1781_),
    .B(_1836_),
    .Y(_1837_));
 sky130_fd_sc_hd__o21ai_1 _6799_ (.A1(_1635_),
    .A2(_1639_),
    .B1(_1696_),
    .Y(_1838_));
 sky130_fd_sc_hd__xnor2_1 _6800_ (.A(_1695_),
    .B(_1838_),
    .Y(_1839_));
 sky130_fd_sc_hd__nand2_1 _6801_ (.A(_1837_),
    .B(_1839_),
    .Y(_1840_));
 sky130_fd_sc_hd__xor2_1 _6802_ (.A(_1692_),
    .B(_1694_),
    .X(_1841_));
 sky130_fd_sc_hd__a21bo_1 _6803_ (.A1(_1733_),
    .A2(_1734_),
    .B1_N(_1780_),
    .X(_1842_));
 sky130_fd_sc_hd__xnor2_1 _6804_ (.A(_1779_),
    .B(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__nand2_1 _6805_ (.A(_1841_),
    .B(_1843_),
    .Y(_1844_));
 sky130_fd_sc_hd__o21ai_1 _6806_ (.A1(_1685_),
    .A2(_1690_),
    .B1(_1641_),
    .Y(_1846_));
 sky130_fd_sc_hd__nor2_1 _6807_ (.A(_1686_),
    .B(_1689_),
    .Y(_1847_));
 sky130_fd_sc_hd__xnor2_1 _6808_ (.A(_1846_),
    .B(_1847_),
    .Y(_1848_));
 sky130_fd_sc_hd__inv_2 _6809_ (.A(_1778_),
    .Y(_1849_));
 sky130_fd_sc_hd__nand2_1 _6810_ (.A(_1735_),
    .B(_1849_),
    .Y(_1850_));
 sky130_fd_sc_hd__nor2_1 _6811_ (.A(_1775_),
    .B(_1777_),
    .Y(_1851_));
 sky130_fd_sc_hd__xnor2_1 _6812_ (.A(_1850_),
    .B(_1851_),
    .Y(_1852_));
 sky130_fd_sc_hd__nor2_1 _6813_ (.A(_1848_),
    .B(_1852_),
    .Y(_1853_));
 sky130_fd_sc_hd__nor2_1 _6814_ (.A(_1642_),
    .B(_1683_),
    .Y(_1854_));
 sky130_fd_sc_hd__xnor2_2 _6815_ (.A(_1688_),
    .B(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__and3_1 _6816_ (.A(_1776_),
    .B(_1738_),
    .C(_1773_),
    .X(_1856_));
 sky130_fd_sc_hd__or2_1 _6817_ (.A(_1777_),
    .B(_1856_),
    .X(_1857_));
 sky130_fd_sc_hd__nor3_1 _6818_ (.A(_1682_),
    .B(_1643_),
    .C(_1680_),
    .Y(_1858_));
 sky130_fd_sc_hd__or2_4 _6819_ (.A(_1683_),
    .B(_1858_),
    .X(_1859_));
 sky130_fd_sc_hd__a211o_1 _6820_ (.A1(_1738_),
    .A2(_1772_),
    .B1(_1739_),
    .C1(_1770_),
    .X(_1860_));
 sky130_fd_sc_hd__nand2_1 _6821_ (.A(_1773_),
    .B(_1860_),
    .Y(_1861_));
 sky130_fd_sc_hd__nor2_1 _6822_ (.A(_1859_),
    .B(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__nor3_1 _6823_ (.A(_1644_),
    .B(_1677_),
    .C(_1679_),
    .Y(_1863_));
 sky130_fd_sc_hd__nor2_1 _6824_ (.A(_1680_),
    .B(_1863_),
    .Y(_1864_));
 sky130_fd_sc_hd__nor3_1 _6825_ (.A(_1740_),
    .B(_1767_),
    .C(_1769_),
    .Y(_1865_));
 sky130_fd_sc_hd__nor2_1 _6826_ (.A(_1770_),
    .B(_1865_),
    .Y(_1867_));
 sky130_fd_sc_hd__and2_1 _6827_ (.A(_1864_),
    .B(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__nor3_1 _6828_ (.A(_1675_),
    .B(_1645_),
    .C(_1673_),
    .Y(_1869_));
 sky130_fd_sc_hd__or2_4 _6829_ (.A(_1677_),
    .B(_1869_),
    .X(_1870_));
 sky130_fd_sc_hd__nor3_1 _6830_ (.A(_1766_),
    .B(_1741_),
    .C(_1764_),
    .Y(_1871_));
 sky130_fd_sc_hd__or2_1 _6831_ (.A(_1767_),
    .B(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__xor2_2 _6832_ (.A(_1870_),
    .B(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__a211oi_1 _6833_ (.A1(_1672_),
    .A2(_1671_),
    .B1(_1670_),
    .C1(_1646_),
    .Y(_1874_));
 sky130_fd_sc_hd__nor2_1 _6834_ (.A(_1673_),
    .B(_1874_),
    .Y(_1875_));
 sky130_fd_sc_hd__a211oi_1 _6835_ (.A1(_1763_),
    .A2(_1762_),
    .B1(_1761_),
    .C1(_1742_),
    .Y(_1876_));
 sky130_fd_sc_hd__nor2_1 _6836_ (.A(_1764_),
    .B(_1876_),
    .Y(_1877_));
 sky130_fd_sc_hd__xor2_1 _6837_ (.A(_1875_),
    .B(_1877_),
    .X(_1878_));
 sky130_fd_sc_hd__a211oi_1 _6838_ (.A1(_1668_),
    .A2(_1669_),
    .B1(_1647_),
    .C1(_1667_),
    .Y(_1879_));
 sky130_fd_sc_hd__or2_1 _6839_ (.A(_1670_),
    .B(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__a211oi_1 _6840_ (.A1(_1759_),
    .A2(_1760_),
    .B1(_1743_),
    .C1(_1758_),
    .Y(_1881_));
 sky130_fd_sc_hd__or2_1 _6841_ (.A(_1761_),
    .B(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__nand2_1 _6842_ (.A(_1880_),
    .B(_1882_),
    .Y(_1883_));
 sky130_fd_sc_hd__and2_1 _6843_ (.A(_1652_),
    .B(_1659_),
    .X(_1884_));
 sky130_fd_sc_hd__xnor2_2 _6844_ (.A(_1661_),
    .B(_1884_),
    .Y(_1885_));
 sky130_fd_sc_hd__nor2_1 _6845_ (.A(_1744_),
    .B(_1746_),
    .Y(_1886_));
 sky130_fd_sc_hd__a22oi_1 _6846_ (.A1(_3576_),
    .A2(\M1.U1.U2.u2.instance11_10.Prop_L ),
    .B1(\In2_reg[2] ),
    .B2(_3426_),
    .Y(_1888_));
 sky130_fd_sc_hd__or2_1 _6847_ (.A(_1745_),
    .B(_1888_),
    .X(_1889_));
 sky130_fd_sc_hd__nor2_2 _6848_ (.A(_1886_),
    .B(_1889_),
    .Y(_1890_));
 sky130_fd_sc_hd__o21a_1 _6849_ (.A1(_1745_),
    .A2(_1890_),
    .B1(_1751_),
    .X(_1891_));
 sky130_fd_sc_hd__nor3_1 _6850_ (.A(_1745_),
    .B(_1751_),
    .C(_1890_),
    .Y(_1892_));
 sky130_fd_sc_hd__or2_1 _6851_ (.A(_1891_),
    .B(_1892_),
    .X(_1893_));
 sky130_fd_sc_hd__xor2_1 _6852_ (.A(_1885_),
    .B(_1893_),
    .X(_1894_));
 sky130_fd_sc_hd__xor2_2 _6853_ (.A(_1658_),
    .B(_1654_),
    .X(_1895_));
 sky130_fd_sc_hd__a22oi_1 _6854_ (.A1(net126),
    .A2(_1617_),
    .B1(_1712_),
    .B2(_3576_),
    .Y(_1896_));
 sky130_fd_sc_hd__nor2_1 _6855_ (.A(_1746_),
    .B(_1896_),
    .Y(_1897_));
 sky130_fd_sc_hd__xnor2_1 _6856_ (.A(_1744_),
    .B(_1897_),
    .Y(_1898_));
 sky130_fd_sc_hd__and2_1 _6857_ (.A(_1895_),
    .B(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__a41o_1 _6858_ (.A1(_3586_),
    .A2(_3503_),
    .A3(_1622_),
    .A4(_1626_),
    .B1(_1656_),
    .X(_1900_));
 sky130_fd_sc_hd__nand4_1 _6859_ (.A(_3437_),
    .B(_3586_),
    .C(_1622_),
    .D(_1626_),
    .Y(_1901_));
 sky130_fd_sc_hd__a22o_1 _6860_ (.A1(_3576_),
    .A2(_1621_),
    .B1(_1626_),
    .B2(_3426_),
    .X(_1902_));
 sky130_fd_sc_hd__nand2_1 _6861_ (.A(_1901_),
    .B(_1902_),
    .Y(_1903_));
 sky130_fd_sc_hd__xnor2_1 _6862_ (.A(_1900_),
    .B(_1903_),
    .Y(_1904_));
 sky130_fd_sc_hd__nand2_1 _6863_ (.A(_3536_),
    .B(_1626_),
    .Y(_1905_));
 sky130_fd_sc_hd__a32o_1 _6864_ (.A1(_3503_),
    .A2(_1622_),
    .A3(_1905_),
    .B1(_1626_),
    .B2(_3586_),
    .X(_1906_));
 sky130_fd_sc_hd__a22oi_1 _6865_ (.A1(_3536_),
    .A2(_1617_),
    .B1(_1712_),
    .B2(net126),
    .Y(_1907_));
 sky130_fd_sc_hd__nor2_1 _6866_ (.A(_1744_),
    .B(_1907_),
    .Y(_1909_));
 sky130_fd_sc_hd__a31o_1 _6867_ (.A1(_3546_),
    .A2(_1712_),
    .A3(_1906_),
    .B1(_1909_),
    .X(_1910_));
 sky130_fd_sc_hd__and4_1 _6868_ (.A(_3546_),
    .B(_1712_),
    .C(_1909_),
    .D(_1906_),
    .X(_1911_));
 sky130_fd_sc_hd__a21oi_1 _6869_ (.A1(_1904_),
    .A2(_1910_),
    .B1(_1911_),
    .Y(_1912_));
 sky130_fd_sc_hd__or2_1 _6870_ (.A(_1895_),
    .B(_1898_),
    .X(_1913_));
 sky130_fd_sc_hd__o21ai_1 _6871_ (.A1(_1899_),
    .A2(_1912_),
    .B1(_1913_),
    .Y(_1914_));
 sky130_fd_sc_hd__a21bo_1 _6872_ (.A1(_1622_),
    .A2(_1650_),
    .B1_N(_1655_),
    .X(_1915_));
 sky130_fd_sc_hd__a21oi_2 _6873_ (.A1(_1658_),
    .A2(_1653_),
    .B1(_1651_),
    .Y(_1916_));
 sky130_fd_sc_hd__xnor2_1 _6874_ (.A(_1916_),
    .B(_1915_),
    .Y(_1917_));
 sky130_fd_sc_hd__nand2_1 _6875_ (.A(_1886_),
    .B(_1889_),
    .Y(_1918_));
 sky130_fd_sc_hd__and2b_1 _6876_ (.A_N(_1890_),
    .B(_1918_),
    .X(_1919_));
 sky130_fd_sc_hd__xnor2_1 _6877_ (.A(_1917_),
    .B(_1919_),
    .Y(_1920_));
 sky130_fd_sc_hd__and2b_1 _6878_ (.A_N(_1917_),
    .B(_1919_),
    .X(_1921_));
 sky130_fd_sc_hd__a21o_1 _6879_ (.A1(_1914_),
    .A2(_1920_),
    .B1(_1921_),
    .X(_1922_));
 sky130_fd_sc_hd__nor2_1 _6880_ (.A(_1885_),
    .B(_1893_),
    .Y(_1923_));
 sky130_fd_sc_hd__a21o_1 _6881_ (.A1(_1894_),
    .A2(_1922_),
    .B1(_1923_),
    .X(_1924_));
 sky130_fd_sc_hd__o21ba_1 _6882_ (.A1(_1661_),
    .A2(_1884_),
    .B1_N(_1648_),
    .X(_1925_));
 sky130_fd_sc_hd__xnor2_2 _6883_ (.A(_1663_),
    .B(_1925_),
    .Y(_1926_));
 sky130_fd_sc_hd__a211o_1 _6884_ (.A1(_1752_),
    .A2(_1754_),
    .B1(_1891_),
    .C1(_1748_),
    .X(_1927_));
 sky130_fd_sc_hd__o211ai_1 _6885_ (.A1(_1748_),
    .A2(_1891_),
    .B1(_1754_),
    .C1(_1752_),
    .Y(_1928_));
 sky130_fd_sc_hd__nand2_1 _6886_ (.A(_1927_),
    .B(_1928_),
    .Y(_1930_));
 sky130_fd_sc_hd__nand2_1 _6887_ (.A(_1926_),
    .B(_1930_),
    .Y(_1931_));
 sky130_fd_sc_hd__nor2_1 _6888_ (.A(_1926_),
    .B(_1930_),
    .Y(_1932_));
 sky130_fd_sc_hd__a21o_1 _6889_ (.A1(_1924_),
    .A2(_1931_),
    .B1(_1932_),
    .X(_1933_));
 sky130_fd_sc_hd__a2111oi_1 _6890_ (.A1(_1666_),
    .A2(_1665_),
    .B1(_1664_),
    .C1(_1649_),
    .D1(_1648_),
    .Y(_1934_));
 sky130_fd_sc_hd__nor2_1 _6891_ (.A(_1667_),
    .B(_1934_),
    .Y(_1935_));
 sky130_fd_sc_hd__a211oi_1 _6892_ (.A1(_1757_),
    .A2(_1756_),
    .B1(_1755_),
    .C1(_1753_),
    .Y(_1936_));
 sky130_fd_sc_hd__nor2_1 _6893_ (.A(_1758_),
    .B(_1936_),
    .Y(_1937_));
 sky130_fd_sc_hd__and2_1 _6894_ (.A(_1935_),
    .B(_1937_),
    .X(_1938_));
 sky130_fd_sc_hd__nor2_1 _6895_ (.A(_1935_),
    .B(_1937_),
    .Y(_1939_));
 sky130_fd_sc_hd__nor2_1 _6896_ (.A(_1938_),
    .B(_1939_),
    .Y(_1940_));
 sky130_fd_sc_hd__nor2_1 _6897_ (.A(_1880_),
    .B(_1882_),
    .Y(_1941_));
 sky130_fd_sc_hd__a211o_1 _6898_ (.A1(_1933_),
    .A2(_1940_),
    .B1(_1941_),
    .C1(_1938_),
    .X(_1942_));
 sky130_fd_sc_hd__and2_1 _6899_ (.A(_1875_),
    .B(_1877_),
    .X(_1943_));
 sky130_fd_sc_hd__a31o_1 _6900_ (.A1(_1878_),
    .A2(_1883_),
    .A3(_1942_),
    .B1(_1943_),
    .X(_1944_));
 sky130_fd_sc_hd__nor2_1 _6901_ (.A(_1870_),
    .B(_1872_),
    .Y(_1945_));
 sky130_fd_sc_hd__a21o_1 _6902_ (.A1(_1873_),
    .A2(_1944_),
    .B1(_1945_),
    .X(_1946_));
 sky130_fd_sc_hd__xor2_1 _6903_ (.A(_1864_),
    .B(_1867_),
    .X(_1947_));
 sky130_fd_sc_hd__and2_1 _6904_ (.A(_1946_),
    .B(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__xor2_1 _6905_ (.A(_1859_),
    .B(_1861_),
    .X(_1949_));
 sky130_fd_sc_hd__o21a_1 _6906_ (.A1(_1868_),
    .A2(_1948_),
    .B1(_1949_),
    .X(_1951_));
 sky130_fd_sc_hd__xor2_1 _6907_ (.A(_1855_),
    .B(_1857_),
    .X(_1952_));
 sky130_fd_sc_hd__o21a_1 _6908_ (.A1(_1862_),
    .A2(_1951_),
    .B1(_1952_),
    .X(_1953_));
 sky130_fd_sc_hd__o21bai_4 _6909_ (.A1(_1855_),
    .A2(_1857_),
    .B1_N(_1953_),
    .Y(_1954_));
 sky130_fd_sc_hd__nand2_1 _6910_ (.A(_1848_),
    .B(_1852_),
    .Y(_1955_));
 sky130_fd_sc_hd__or2_1 _6911_ (.A(_1841_),
    .B(_1843_),
    .X(_1956_));
 sky130_fd_sc_hd__and2_4 _6912_ (.A(_1844_),
    .B(_1956_),
    .X(_1957_));
 sky130_fd_sc_hd__o211ai_2 _6913_ (.A1(_1853_),
    .A2(_1954_),
    .B1(_1955_),
    .C1(_1957_),
    .Y(_1958_));
 sky130_fd_sc_hd__or2_1 _6914_ (.A(_1837_),
    .B(_1839_),
    .X(_1959_));
 sky130_fd_sc_hd__inv_2 _6915_ (.A(_1959_),
    .Y(_1960_));
 sky130_fd_sc_hd__xnor2_1 _6916_ (.A(_1832_),
    .B(_1835_),
    .Y(_1961_));
 sky130_fd_sc_hd__a311oi_2 _6917_ (.A1(_1840_),
    .A2(_1844_),
    .A3(_1958_),
    .B1(_1960_),
    .C1(_1961_),
    .Y(_1962_));
 sky130_fd_sc_hd__a21o_1 _6918_ (.A1(_1832_),
    .A2(_1835_),
    .B1(_1962_),
    .X(_1963_));
 sky130_fd_sc_hd__nand2b_1 _6919_ (.A_N(_1830_),
    .B(_1828_),
    .Y(_1964_));
 sky130_fd_sc_hd__xor2_1 _6920_ (.A(_1822_),
    .B(_1825_),
    .X(_1965_));
 sky130_fd_sc_hd__o211a_1 _6921_ (.A1(_1831_),
    .A2(_1963_),
    .B1(_1964_),
    .C1(_1965_),
    .X(_1966_));
 sky130_fd_sc_hd__nor2_1 _6922_ (.A(_1705_),
    .B(_1817_),
    .Y(_1967_));
 sky130_fd_sc_hd__xnor2_1 _6923_ (.A(_1967_),
    .B(_1819_),
    .Y(_1968_));
 sky130_fd_sc_hd__o21ai_1 _6924_ (.A1(_1826_),
    .A2(_1966_),
    .B1(_1968_),
    .Y(_1969_));
 sky130_fd_sc_hd__nor2b_4 _6925_ (.A(_1709_),
    .B_N(_1815_),
    .Y(_1970_));
 sky130_fd_sc_hd__xnor2_2 _6926_ (.A(_1814_),
    .B(_1970_),
    .Y(_1972_));
 sky130_fd_sc_hd__a21bo_1 _6927_ (.A1(_1820_),
    .A2(_1969_),
    .B1_N(_1972_),
    .X(_1973_));
 sky130_fd_sc_hd__xor2_1 _6928_ (.A(_1806_),
    .B(_1810_),
    .X(_1974_));
 sky130_fd_sc_hd__a21o_1 _6929_ (.A1(_1973_),
    .A2(_1816_),
    .B1(_1974_),
    .X(_1975_));
 sky130_fd_sc_hd__a21oi_1 _6930_ (.A1(_1625_),
    .A2(_1801_),
    .B1(_1802_),
    .Y(_1976_));
 sky130_fd_sc_hd__or2_4 _6931_ (.A(_1803_),
    .B(_1976_),
    .X(_1977_));
 sky130_fd_sc_hd__a21oi_2 _6932_ (.A1(_1811_),
    .A2(_1975_),
    .B1(_1977_),
    .Y(_1978_));
 sky130_fd_sc_hd__xnor2_1 _6933_ (.A(_1801_),
    .B(_1800_),
    .Y(_1979_));
 sky130_fd_sc_hd__o21ai_1 _6934_ (.A1(_1803_),
    .A2(_1978_),
    .B1(_1979_),
    .Y(_1980_));
 sky130_fd_sc_hd__a21bo_2 _6935_ (.A1(_1711_),
    .A2(_1800_),
    .B1_N(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__nor2_1 _6936_ (.A(_1799_),
    .B(_1716_),
    .Y(_1982_));
 sky130_fd_sc_hd__a21bo_1 _6937_ (.A1(_1620_),
    .A2(_1981_),
    .B1_N(_1982_),
    .X(_1983_));
 sky130_fd_sc_hd__nor3_1 _6938_ (.A(_1603_),
    .B(_1447_),
    .C(_1602_),
    .Y(_1984_));
 sky130_fd_sc_hd__or2_1 _6939_ (.A(_1604_),
    .B(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__xnor2_2 _6940_ (.A(_1983_),
    .B(_1985_),
    .Y(_1986_));
 sky130_fd_sc_hd__nand2_1 _6941_ (.A(_1620_),
    .B(_1982_),
    .Y(_1987_));
 sky130_fd_sc_hd__xor2_2 _6942_ (.A(_1981_),
    .B(_1987_),
    .X(_1988_));
 sky130_fd_sc_hd__nor3_1 _6943_ (.A(_1601_),
    .B(_1452_),
    .C(_1600_),
    .Y(_1989_));
 sky130_fd_sc_hd__or2_1 _6944_ (.A(_1602_),
    .B(_1989_),
    .X(_1990_));
 sky130_fd_sc_hd__xnor2_2 _6945_ (.A(_1988_),
    .B(_1990_),
    .Y(_1991_));
 sky130_fd_sc_hd__or3_4 _6946_ (.A(_1979_),
    .B(_1803_),
    .C(_1978_),
    .X(_1993_));
 sky130_fd_sc_hd__nand2_4 _6947_ (.A(_1980_),
    .B(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__nor2_1 _6948_ (.A(_1455_),
    .B(_1598_),
    .Y(_1995_));
 sky130_fd_sc_hd__xnor2_1 _6949_ (.A(_1599_),
    .B(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__xor2_4 _6950_ (.A(_1994_),
    .B(_1996_),
    .X(_1997_));
 sky130_fd_sc_hd__and3_1 _6951_ (.A(_1977_),
    .B(_1811_),
    .C(_1975_),
    .X(_1998_));
 sky130_fd_sc_hd__or2_4 _6952_ (.A(_1978_),
    .B(_1998_),
    .X(_1999_));
 sky130_fd_sc_hd__and3_1 _6953_ (.A(_1597_),
    .B(_1462_),
    .C(_1595_),
    .X(_2000_));
 sky130_fd_sc_hd__or2_1 _6954_ (.A(_1598_),
    .B(_2000_),
    .X(_2001_));
 sky130_fd_sc_hd__xor2_2 _6955_ (.A(_1999_),
    .B(_2001_),
    .X(_2002_));
 sky130_fd_sc_hd__nand3_1 _6956_ (.A(_1816_),
    .B(_1973_),
    .C(_1974_),
    .Y(_2003_));
 sky130_fd_sc_hd__nand2_1 _6957_ (.A(_1975_),
    .B(_2003_),
    .Y(_2004_));
 sky130_fd_sc_hd__nand3_1 _6958_ (.A(_1465_),
    .B(_1593_),
    .C(_1594_),
    .Y(_2005_));
 sky130_fd_sc_hd__nand2_1 _6959_ (.A(_1595_),
    .B(_2005_),
    .Y(_2006_));
 sky130_fd_sc_hd__nand2_1 _6960_ (.A(_2004_),
    .B(_2006_),
    .Y(_2007_));
 sky130_fd_sc_hd__o21ai_1 _6961_ (.A1(_1831_),
    .A2(_1963_),
    .B1(_1964_),
    .Y(_2008_));
 sky130_fd_sc_hd__xnor2_1 _6962_ (.A(_1965_),
    .B(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__nor3_1 _6963_ (.A(_1586_),
    .B(_1479_),
    .C(_1584_),
    .Y(_2010_));
 sky130_fd_sc_hd__nor2_1 _6964_ (.A(_1587_),
    .B(_2010_),
    .Y(_2011_));
 sky130_fd_sc_hd__and2_1 _6965_ (.A(_2009_),
    .B(_2011_),
    .X(_2012_));
 sky130_fd_sc_hd__nor2_1 _6966_ (.A(_2009_),
    .B(_2011_),
    .Y(_2014_));
 sky130_fd_sc_hd__nor2_1 _6967_ (.A(_2012_),
    .B(_2014_),
    .Y(_2015_));
 sky130_fd_sc_hd__and3_1 _6968_ (.A(_1583_),
    .B(_1483_),
    .C(_1581_),
    .X(_2016_));
 sky130_fd_sc_hd__or2_1 _6969_ (.A(_1584_),
    .B(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__nor2b_1 _6970_ (.A(_1831_),
    .B_N(_1964_),
    .Y(_2018_));
 sky130_fd_sc_hd__xnor2_1 _6971_ (.A(_1963_),
    .B(_2018_),
    .Y(_2019_));
 sky130_fd_sc_hd__nand2_1 _6972_ (.A(_2017_),
    .B(_2019_),
    .Y(_2020_));
 sky130_fd_sc_hd__and2_4 _6973_ (.A(_1844_),
    .B(_1958_),
    .X(_2021_));
 sky130_fd_sc_hd__o211a_1 _6974_ (.A1(_1960_),
    .A2(_2021_),
    .B1(_1840_),
    .C1(_1961_),
    .X(_2022_));
 sky130_fd_sc_hd__nor2_1 _6975_ (.A(_1962_),
    .B(_2022_),
    .Y(_2023_));
 sky130_fd_sc_hd__or3_1 _6976_ (.A(_1580_),
    .B(_1488_),
    .C(_1579_),
    .X(_2024_));
 sky130_fd_sc_hd__and2_1 _6977_ (.A(_1581_),
    .B(_2024_),
    .X(_2025_));
 sky130_fd_sc_hd__xor2_2 _6978_ (.A(_2023_),
    .B(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__nor2_1 _6979_ (.A(_1492_),
    .B(_1576_),
    .Y(_2027_));
 sky130_fd_sc_hd__xnor2_2 _6980_ (.A(_1578_),
    .B(_2027_),
    .Y(_2028_));
 sky130_fd_sc_hd__nand2_1 _6981_ (.A(_1959_),
    .B(_1840_),
    .Y(_2029_));
 sky130_fd_sc_hd__xnor2_2 _6982_ (.A(_2021_),
    .B(_2029_),
    .Y(_2030_));
 sky130_fd_sc_hd__xor2_2 _6983_ (.A(_2028_),
    .B(_2030_),
    .X(_2031_));
 sky130_fd_sc_hd__o21ai_2 _6984_ (.A1(_1853_),
    .A2(_1954_),
    .B1(_1955_),
    .Y(_2032_));
 sky130_fd_sc_hd__xnor2_2 _6985_ (.A(_2032_),
    .B(_1957_),
    .Y(_2033_));
 sky130_fd_sc_hd__nor3_1 _6986_ (.A(_1500_),
    .B(_1573_),
    .C(_1575_),
    .Y(_2035_));
 sky130_fd_sc_hd__nor2_1 _6987_ (.A(_1576_),
    .B(_2035_),
    .Y(_2036_));
 sky130_fd_sc_hd__xor2_2 _6988_ (.A(_2033_),
    .B(_2036_),
    .X(_2037_));
 sky130_fd_sc_hd__nor3_1 _6989_ (.A(_1572_),
    .B(_1504_),
    .C(_1571_),
    .Y(_2038_));
 sky130_fd_sc_hd__or2_1 _6990_ (.A(_1573_),
    .B(_2038_),
    .X(_2039_));
 sky130_fd_sc_hd__and2b_1 _6991_ (.A_N(_1853_),
    .B(_1955_),
    .X(_2040_));
 sky130_fd_sc_hd__xnor2_2 _6992_ (.A(_2040_),
    .B(_1954_),
    .Y(_2041_));
 sky130_fd_sc_hd__xor2_1 _6993_ (.A(_2039_),
    .B(_2041_),
    .X(_2042_));
 sky130_fd_sc_hd__nor3_1 _6994_ (.A(_1570_),
    .B(_1509_),
    .C(_1568_),
    .Y(_2043_));
 sky130_fd_sc_hd__nor2_1 _6995_ (.A(_1571_),
    .B(_2043_),
    .Y(_2044_));
 sky130_fd_sc_hd__nor3_1 _6996_ (.A(_1952_),
    .B(_1862_),
    .C(_1951_),
    .Y(_2045_));
 sky130_fd_sc_hd__nor2_1 _6997_ (.A(_1953_),
    .B(_2045_),
    .Y(_2046_));
 sky130_fd_sc_hd__xor2_1 _6998_ (.A(_2044_),
    .B(_2046_),
    .X(_2047_));
 sky130_fd_sc_hd__nor3_1 _6999_ (.A(_1949_),
    .B(_1868_),
    .C(_1948_),
    .Y(_2048_));
 sky130_fd_sc_hd__nor2_1 _7000_ (.A(_1951_),
    .B(_2048_),
    .Y(_2049_));
 sky130_fd_sc_hd__nor3_1 _7001_ (.A(_1567_),
    .B(_1512_),
    .C(_1565_),
    .Y(_2050_));
 sky130_fd_sc_hd__nor2_1 _7002_ (.A(_1568_),
    .B(_2050_),
    .Y(_2051_));
 sky130_fd_sc_hd__xor2_1 _7003_ (.A(_2049_),
    .B(_2051_),
    .X(_2052_));
 sky130_fd_sc_hd__nor3_1 _7004_ (.A(_1564_),
    .B(_1517_),
    .C(_1562_),
    .Y(_2053_));
 sky130_fd_sc_hd__or2_1 _7005_ (.A(_1565_),
    .B(_2053_),
    .X(_2054_));
 sky130_fd_sc_hd__inv_2 _7006_ (.A(_2054_),
    .Y(_2056_));
 sky130_fd_sc_hd__nor2_1 _7007_ (.A(_1946_),
    .B(_1947_),
    .Y(_2057_));
 sky130_fd_sc_hd__nor2_1 _7008_ (.A(_1948_),
    .B(_2057_),
    .Y(_2058_));
 sky130_fd_sc_hd__nor2_1 _7009_ (.A(_2056_),
    .B(_2058_),
    .Y(_2059_));
 sky130_fd_sc_hd__nor3_1 _7010_ (.A(_1561_),
    .B(_1522_),
    .C(_1559_),
    .Y(_2060_));
 sky130_fd_sc_hd__nor2_1 _7011_ (.A(_1562_),
    .B(_2060_),
    .Y(_2061_));
 sky130_fd_sc_hd__xnor2_2 _7012_ (.A(_1873_),
    .B(_1944_),
    .Y(_2062_));
 sky130_fd_sc_hd__xor2_1 _7013_ (.A(_2061_),
    .B(_2062_),
    .X(_2063_));
 sky130_fd_sc_hd__inv_2 _7014_ (.A(_2063_),
    .Y(_2064_));
 sky130_fd_sc_hd__nand2_1 _7015_ (.A(_1883_),
    .B(_1942_),
    .Y(_2065_));
 sky130_fd_sc_hd__xnor2_1 _7016_ (.A(_1878_),
    .B(_2065_),
    .Y(_2067_));
 sky130_fd_sc_hd__or2_1 _7017_ (.A(_1527_),
    .B(_1556_),
    .X(_2068_));
 sky130_fd_sc_hd__xnor2_1 _7018_ (.A(_1558_),
    .B(_2068_),
    .Y(_2069_));
 sky130_fd_sc_hd__xnor2_1 _7019_ (.A(_2067_),
    .B(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__nor3_1 _7020_ (.A(_1555_),
    .B(_1535_),
    .C(_1553_),
    .Y(_2071_));
 sky130_fd_sc_hd__nor2_1 _7021_ (.A(_1556_),
    .B(_2071_),
    .Y(_2072_));
 sky130_fd_sc_hd__a21o_1 _7022_ (.A1(_1933_),
    .A2(_1940_),
    .B1(_1938_),
    .X(_2073_));
 sky130_fd_sc_hd__nand2b_1 _7023_ (.A_N(_1941_),
    .B(_1883_),
    .Y(_2074_));
 sky130_fd_sc_hd__xnor2_1 _7024_ (.A(_2073_),
    .B(_2074_),
    .Y(_2075_));
 sky130_fd_sc_hd__xnor2_1 _7025_ (.A(_2072_),
    .B(_2075_),
    .Y(_2076_));
 sky130_fd_sc_hd__xor2_2 _7026_ (.A(_1933_),
    .B(_1940_),
    .X(_2077_));
 sky130_fd_sc_hd__nor3_1 _7027_ (.A(_1552_),
    .B(_1541_),
    .C(_1550_),
    .Y(_2078_));
 sky130_fd_sc_hd__nor2_1 _7028_ (.A(_1553_),
    .B(_2078_),
    .Y(_2079_));
 sky130_fd_sc_hd__xnor2_1 _7029_ (.A(_2077_),
    .B(_2079_),
    .Y(_2080_));
 sky130_fd_sc_hd__xnor2_1 _7030_ (.A(_1926_),
    .B(_1930_),
    .Y(_2081_));
 sky130_fd_sc_hd__xnor2_1 _7031_ (.A(_1924_),
    .B(_2081_),
    .Y(_2082_));
 sky130_fd_sc_hd__xnor2_1 _7032_ (.A(_1543_),
    .B(_1549_),
    .Y(_2083_));
 sky130_fd_sc_hd__nand2_1 _7033_ (.A(_2082_),
    .B(_2083_),
    .Y(_2084_));
 sky130_fd_sc_hd__xor2_1 _7034_ (.A(_1894_),
    .B(_1922_),
    .X(_2085_));
 sky130_fd_sc_hd__nand2_1 _7035_ (.A(_1914_),
    .B(_1920_),
    .Y(_2086_));
 sky130_fd_sc_hd__xor2_1 _7036_ (.A(_1895_),
    .B(_1898_),
    .X(_2088_));
 sky130_fd_sc_hd__xnor2_1 _7037_ (.A(_2088_),
    .B(_1912_),
    .Y(_2089_));
 sky130_fd_sc_hd__a22oi_1 _7038_ (.A1(_3556_),
    .A2(_1348_),
    .B1(_1353_),
    .B2(_3525_),
    .Y(_2090_));
 sky130_fd_sc_hd__nor2_1 _7039_ (.A(_1394_),
    .B(_2090_),
    .Y(_2091_));
 sky130_fd_sc_hd__a21o_1 _7040_ (.A1(_1546_),
    .A2(_2089_),
    .B1(_2091_),
    .X(_2092_));
 sky130_fd_sc_hd__or2_1 _7041_ (.A(_1914_),
    .B(_1920_),
    .X(_2093_));
 sky130_fd_sc_hd__and3_1 _7042_ (.A(_1546_),
    .B(_2091_),
    .C(_2089_),
    .X(_2094_));
 sky130_fd_sc_hd__a31o_1 _7043_ (.A1(_2086_),
    .A2(_2092_),
    .A3(_2093_),
    .B1(_2094_),
    .X(_2095_));
 sky130_fd_sc_hd__nand2_1 _7044_ (.A(_2085_),
    .B(_2095_),
    .Y(_2096_));
 sky130_fd_sc_hd__nor2_1 _7045_ (.A(_2085_),
    .B(_2095_),
    .Y(_2097_));
 sky130_fd_sc_hd__a21oi_1 _7046_ (.A1(_3556_),
    .A2(_1256_),
    .B1(_1548_),
    .Y(_2098_));
 sky130_fd_sc_hd__or3_1 _7047_ (.A(_1549_),
    .B(_2097_),
    .C(_2098_),
    .X(_2099_));
 sky130_fd_sc_hd__nor2_1 _7048_ (.A(_2082_),
    .B(_2083_),
    .Y(_2100_));
 sky130_fd_sc_hd__a31o_1 _7049_ (.A1(_2084_),
    .A2(_2096_),
    .A3(_2099_),
    .B1(_2100_),
    .X(_2101_));
 sky130_fd_sc_hd__nand2_1 _7050_ (.A(_2077_),
    .B(_2079_),
    .Y(_2102_));
 sky130_fd_sc_hd__o21a_1 _7051_ (.A1(_2080_),
    .A2(_2101_),
    .B1(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__nand2_1 _7052_ (.A(_2072_),
    .B(_2075_),
    .Y(_2104_));
 sky130_fd_sc_hd__o21ai_1 _7053_ (.A1(_2076_),
    .A2(_2103_),
    .B1(_2104_),
    .Y(_2105_));
 sky130_fd_sc_hd__inv_2 _7054_ (.A(_2069_),
    .Y(_2106_));
 sky130_fd_sc_hd__and2_1 _7055_ (.A(_2067_),
    .B(_2106_),
    .X(_2107_));
 sky130_fd_sc_hd__a21o_1 _7056_ (.A1(_2070_),
    .A2(_2105_),
    .B1(_2107_),
    .X(_2109_));
 sky130_fd_sc_hd__inv_2 _7057_ (.A(_2061_),
    .Y(_2110_));
 sky130_fd_sc_hd__nor2_1 _7058_ (.A(_2110_),
    .B(_2062_),
    .Y(_2111_));
 sky130_fd_sc_hd__a21oi_1 _7059_ (.A1(_2064_),
    .A2(_2109_),
    .B1(_2111_),
    .Y(_2112_));
 sky130_fd_sc_hd__and2_1 _7060_ (.A(_2056_),
    .B(_2058_),
    .X(_2113_));
 sky130_fd_sc_hd__o21bai_1 _7061_ (.A1(_2059_),
    .A2(_2112_),
    .B1_N(_2113_),
    .Y(_2114_));
 sky130_fd_sc_hd__and2_1 _7062_ (.A(_2049_),
    .B(_2051_),
    .X(_2115_));
 sky130_fd_sc_hd__a21o_1 _7063_ (.A1(_2052_),
    .A2(_2114_),
    .B1(_2115_),
    .X(_2116_));
 sky130_fd_sc_hd__and2_1 _7064_ (.A(_2044_),
    .B(_2046_),
    .X(_2117_));
 sky130_fd_sc_hd__a21o_1 _7065_ (.A1(_2047_),
    .A2(_2116_),
    .B1(_2117_),
    .X(_2118_));
 sky130_fd_sc_hd__nor2_1 _7066_ (.A(_2039_),
    .B(_2041_),
    .Y(_2119_));
 sky130_fd_sc_hd__a21o_1 _7067_ (.A1(_2118_),
    .A2(_2042_),
    .B1(_2119_),
    .X(_2120_));
 sky130_fd_sc_hd__and2_1 _7068_ (.A(_2033_),
    .B(_2036_),
    .X(_2121_));
 sky130_fd_sc_hd__a21o_1 _7069_ (.A1(_2120_),
    .A2(_2037_),
    .B1(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__nor2_1 _7070_ (.A(_2028_),
    .B(_2030_),
    .Y(_2123_));
 sky130_fd_sc_hd__a21o_1 _7071_ (.A1(_2122_),
    .A2(_2031_),
    .B1(_2123_),
    .X(_2124_));
 sky130_fd_sc_hd__and2_1 _7072_ (.A(_2023_),
    .B(_2025_),
    .X(_2125_));
 sky130_fd_sc_hd__a21o_1 _7073_ (.A1(_2124_),
    .A2(_2026_),
    .B1(_2125_),
    .X(_2126_));
 sky130_fd_sc_hd__nor2_1 _7074_ (.A(_2017_),
    .B(_2019_),
    .Y(_2127_));
 sky130_fd_sc_hd__a21o_1 _7075_ (.A1(_2126_),
    .A2(_2020_),
    .B1(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__a21o_1 _7076_ (.A1(_2128_),
    .A2(_2015_),
    .B1(_2012_),
    .X(_2130_));
 sky130_fd_sc_hd__or3_1 _7077_ (.A(_1968_),
    .B(_1826_),
    .C(_1966_),
    .X(_2131_));
 sky130_fd_sc_hd__nand2_1 _7078_ (.A(_1969_),
    .B(_2131_),
    .Y(_2132_));
 sky130_fd_sc_hd__nor3_1 _7079_ (.A(_1589_),
    .B(_1473_),
    .C(_1587_),
    .Y(_2133_));
 sky130_fd_sc_hd__or2_1 _7080_ (.A(_1590_),
    .B(_2133_),
    .X(_2134_));
 sky130_fd_sc_hd__nor2_1 _7081_ (.A(_2132_),
    .B(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__and2_1 _7082_ (.A(_2132_),
    .B(_2134_),
    .X(_2136_));
 sky130_fd_sc_hd__nor2_1 _7083_ (.A(_2135_),
    .B(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__a21o_4 _7084_ (.A1(_2130_),
    .A2(_2137_),
    .B1(_2135_),
    .X(_2138_));
 sky130_fd_sc_hd__nand3b_1 _7085_ (.A_N(_1972_),
    .B(_1820_),
    .C(_1969_),
    .Y(_2139_));
 sky130_fd_sc_hd__and2_1 _7086_ (.A(_1973_),
    .B(_2139_),
    .X(_2140_));
 sky130_fd_sc_hd__or3_1 _7087_ (.A(_1592_),
    .B(_1470_),
    .C(_1590_),
    .X(_2141_));
 sky130_fd_sc_hd__and2_1 _7088_ (.A(_1593_),
    .B(_2141_),
    .X(_2142_));
 sky130_fd_sc_hd__and2_4 _7089_ (.A(_2140_),
    .B(_2142_),
    .X(_2143_));
 sky130_fd_sc_hd__nor2_2 _7090_ (.A(_2140_),
    .B(_2142_),
    .Y(_2144_));
 sky130_fd_sc_hd__nor2_4 _7091_ (.A(_2144_),
    .B(_2143_),
    .Y(_2145_));
 sky130_fd_sc_hd__nor2_1 _7092_ (.A(_2004_),
    .B(_2006_),
    .Y(_2146_));
 sky130_fd_sc_hd__a211o_4 _7093_ (.A1(_2138_),
    .A2(_2145_),
    .B1(_2146_),
    .C1(_2143_),
    .X(_2147_));
 sky130_fd_sc_hd__nor2_1 _7094_ (.A(_1999_),
    .B(_2001_),
    .Y(_2148_));
 sky130_fd_sc_hd__a31o_4 _7095_ (.A1(_2002_),
    .A2(_2007_),
    .A3(_2147_),
    .B1(_2148_),
    .X(_2149_));
 sky130_fd_sc_hd__nor2_1 _7096_ (.A(_1994_),
    .B(_1996_),
    .Y(_2151_));
 sky130_fd_sc_hd__a21oi_4 _7097_ (.A1(_2149_),
    .A2(_1997_),
    .B1(_2151_),
    .Y(_2152_));
 sky130_fd_sc_hd__or2_1 _7098_ (.A(_1988_),
    .B(_1990_),
    .X(_2153_));
 sky130_fd_sc_hd__o21ai_2 _7099_ (.A1(_2152_),
    .A2(_1991_),
    .B1(_2153_),
    .Y(_2154_));
 sky130_fd_sc_hd__and2b_1 _7100_ (.A_N(_1985_),
    .B(_1983_),
    .X(_2155_));
 sky130_fd_sc_hd__a21oi_2 _7101_ (.A1(_2154_),
    .A2(_1986_),
    .B1(_2155_),
    .Y(_2156_));
 sky130_fd_sc_hd__or3_4 _7102_ (.A(_1613_),
    .B(_1616_),
    .C(_2156_),
    .X(_2157_));
 sky130_fd_sc_hd__xnor2_1 _7103_ (.A(_1346_),
    .B(_1610_),
    .Y(_2158_));
 sky130_fd_sc_hd__nor2_1 _7104_ (.A(_2157_),
    .B(_2158_),
    .Y(_2159_));
 sky130_fd_sc_hd__inv_2 _7105_ (.A(_2159_),
    .Y(_2160_));
 sky130_fd_sc_hd__nor2_1 _7106_ (.A(_1108_),
    .B(_1234_),
    .Y(_2161_));
 sky130_fd_sc_hd__nand2_1 _7107_ (.A(_1235_),
    .B(_2161_),
    .Y(_2162_));
 sky130_fd_sc_hd__or2b_1 _7108_ (.A(_1236_),
    .B_N(_2162_),
    .X(_2163_));
 sky130_fd_sc_hd__a31oi_2 _7109_ (.A1(_1345_),
    .A2(_1611_),
    .A3(_2160_),
    .B1(_2163_),
    .Y(_2164_));
 sky130_fd_sc_hd__o21ai_1 _7110_ (.A1(_1616_),
    .A2(_2156_),
    .B1(_1613_),
    .Y(_2165_));
 sky130_fd_sc_hd__and2_1 _7111_ (.A(_2157_),
    .B(_2165_),
    .X(_2166_));
 sky130_fd_sc_hd__nand3_1 _7112_ (.A(_1231_),
    .B(_1118_),
    .C(_1230_),
    .Y(_2167_));
 sky130_fd_sc_hd__and2_1 _7113_ (.A(_1232_),
    .B(_2167_),
    .X(_2168_));
 sky130_fd_sc_hd__or2_1 _7114_ (.A(_2166_),
    .B(_2168_),
    .X(_2169_));
 sky130_fd_sc_hd__xnor2_1 _7115_ (.A(_1616_),
    .B(_2156_),
    .Y(_2170_));
 sky130_fd_sc_hd__or3_1 _7116_ (.A(_1229_),
    .B(_1123_),
    .C(_1228_),
    .X(_2172_));
 sky130_fd_sc_hd__nand2_1 _7117_ (.A(_1230_),
    .B(_2172_),
    .Y(_2173_));
 sky130_fd_sc_hd__nor2_1 _7118_ (.A(_2170_),
    .B(_2173_),
    .Y(_2174_));
 sky130_fd_sc_hd__and2_1 _7119_ (.A(_2170_),
    .B(_2173_),
    .X(_2175_));
 sky130_fd_sc_hd__nor2_1 _7120_ (.A(_2174_),
    .B(_2175_),
    .Y(_2176_));
 sky130_fd_sc_hd__xnor2_1 _7121_ (.A(_1986_),
    .B(_2154_),
    .Y(_2177_));
 sky130_fd_sc_hd__and3_1 _7122_ (.A(_1227_),
    .B(_1127_),
    .C(_1226_),
    .X(_2178_));
 sky130_fd_sc_hd__or2_1 _7123_ (.A(_1228_),
    .B(_2178_),
    .X(_2179_));
 sky130_fd_sc_hd__nor2_1 _7124_ (.A(_2177_),
    .B(_2179_),
    .Y(_2180_));
 sky130_fd_sc_hd__and2_1 _7125_ (.A(_2177_),
    .B(_2179_),
    .X(_2181_));
 sky130_fd_sc_hd__nor2_1 _7126_ (.A(_2180_),
    .B(_2181_),
    .Y(_2182_));
 sky130_fd_sc_hd__xnor2_2 _7127_ (.A(_1991_),
    .B(_2152_),
    .Y(_2183_));
 sky130_fd_sc_hd__or3_1 _7128_ (.A(_1225_),
    .B(_1132_),
    .C(_1223_),
    .X(_2184_));
 sky130_fd_sc_hd__and2_1 _7129_ (.A(_1226_),
    .B(_2184_),
    .X(_2185_));
 sky130_fd_sc_hd__xnor2_2 _7130_ (.A(_2183_),
    .B(_2185_),
    .Y(_2186_));
 sky130_fd_sc_hd__nand3_1 _7131_ (.A(_1146_),
    .B(_1217_),
    .C(_1218_),
    .Y(_2187_));
 sky130_fd_sc_hd__nand2_1 _7132_ (.A(_1219_),
    .B(_2187_),
    .Y(_2188_));
 sky130_fd_sc_hd__a21o_1 _7133_ (.A1(_2145_),
    .A2(_2138_),
    .B1(_2143_),
    .X(_2189_));
 sky130_fd_sc_hd__and2b_1 _7134_ (.A_N(_2146_),
    .B(_2007_),
    .X(_2190_));
 sky130_fd_sc_hd__xnor2_2 _7135_ (.A(_2189_),
    .B(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hd__xnor2_2 _7136_ (.A(_2191_),
    .B(_2188_),
    .Y(_2193_));
 sky130_fd_sc_hd__xnor2_4 _7137_ (.A(_2138_),
    .B(_2145_),
    .Y(_2194_));
 sky130_fd_sc_hd__nand3_1 _7138_ (.A(_1216_),
    .B(_1151_),
    .C(_1215_),
    .Y(_2195_));
 sky130_fd_sc_hd__nand2_1 _7139_ (.A(_1217_),
    .B(_2195_),
    .Y(_2196_));
 sky130_fd_sc_hd__xor2_2 _7140_ (.A(_2194_),
    .B(_2196_),
    .X(_2197_));
 sky130_fd_sc_hd__nand3_1 _7141_ (.A(_1214_),
    .B(_1155_),
    .C(_1213_),
    .Y(_2198_));
 sky130_fd_sc_hd__nand2_1 _7142_ (.A(_1215_),
    .B(_2198_),
    .Y(_2199_));
 sky130_fd_sc_hd__xnor2_2 _7143_ (.A(_2130_),
    .B(_2137_),
    .Y(_2200_));
 sky130_fd_sc_hd__xor2_1 _7144_ (.A(_2199_),
    .B(_2200_),
    .X(_2201_));
 sky130_fd_sc_hd__xnor2_2 _7145_ (.A(_2015_),
    .B(_2128_),
    .Y(_2202_));
 sky130_fd_sc_hd__or3_1 _7146_ (.A(_1212_),
    .B(_1160_),
    .C(_1210_),
    .X(_2203_));
 sky130_fd_sc_hd__and2_1 _7147_ (.A(_1213_),
    .B(_2203_),
    .X(_2204_));
 sky130_fd_sc_hd__xnor2_1 _7148_ (.A(_2202_),
    .B(_2204_),
    .Y(_2205_));
 sky130_fd_sc_hd__nand2b_1 _7149_ (.A_N(_2127_),
    .B(_2020_),
    .Y(_2206_));
 sky130_fd_sc_hd__xnor2_2 _7150_ (.A(_2206_),
    .B(_2126_),
    .Y(_2207_));
 sky130_fd_sc_hd__and3b_1 _7151_ (.A_N(_1209_),
    .B(_1165_),
    .C(_1208_),
    .X(_2208_));
 sky130_fd_sc_hd__nor2_1 _7152_ (.A(_1210_),
    .B(_2208_),
    .Y(_2209_));
 sky130_fd_sc_hd__xor2_1 _7153_ (.A(_2207_),
    .B(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__xnor2_2 _7154_ (.A(_2026_),
    .B(_2124_),
    .Y(_2211_));
 sky130_fd_sc_hd__nand3_1 _7155_ (.A(_1207_),
    .B(_1170_),
    .C(_1206_),
    .Y(_2212_));
 sky130_fd_sc_hd__nand2_1 _7156_ (.A(_1208_),
    .B(_2212_),
    .Y(_2214_));
 sky130_fd_sc_hd__xor2_1 _7157_ (.A(_2211_),
    .B(_2214_),
    .X(_2215_));
 sky130_fd_sc_hd__xor2_2 _7158_ (.A(_2031_),
    .B(_2122_),
    .X(_2216_));
 sky130_fd_sc_hd__nand3_1 _7159_ (.A(_1205_),
    .B(_1174_),
    .C(_1203_),
    .Y(_2217_));
 sky130_fd_sc_hd__nand2_1 _7160_ (.A(_1206_),
    .B(_2217_),
    .Y(_2218_));
 sky130_fd_sc_hd__xnor2_1 _7161_ (.A(_2216_),
    .B(_2218_),
    .Y(_2219_));
 sky130_fd_sc_hd__xnor2_2 _7162_ (.A(_2037_),
    .B(_2120_),
    .Y(_2220_));
 sky130_fd_sc_hd__or3_1 _7163_ (.A(_1202_),
    .B(_1179_),
    .C(_1200_),
    .X(_2221_));
 sky130_fd_sc_hd__nand2_1 _7164_ (.A(_1203_),
    .B(_2221_),
    .Y(_2222_));
 sky130_fd_sc_hd__xor2_1 _7165_ (.A(_2220_),
    .B(_2222_),
    .X(_2223_));
 sky130_fd_sc_hd__xnor2_1 _7166_ (.A(_2042_),
    .B(_2118_),
    .Y(_2224_));
 sky130_fd_sc_hd__nor3_1 _7167_ (.A(_1183_),
    .B(_1197_),
    .C(_1199_),
    .Y(_2225_));
 sky130_fd_sc_hd__or2_1 _7168_ (.A(_1200_),
    .B(_2225_),
    .X(_2226_));
 sky130_fd_sc_hd__or2_1 _7169_ (.A(_2224_),
    .B(_2226_),
    .X(_2227_));
 sky130_fd_sc_hd__xnor2_1 _7170_ (.A(_2047_),
    .B(_2116_),
    .Y(_2228_));
 sky130_fd_sc_hd__xnor2_1 _7171_ (.A(_1185_),
    .B(_1196_),
    .Y(_2229_));
 sky130_fd_sc_hd__or2_1 _7172_ (.A(_2228_),
    .B(_2229_),
    .X(_2230_));
 sky130_fd_sc_hd__nor2_1 _7173_ (.A(_2113_),
    .B(_2059_),
    .Y(_2231_));
 sky130_fd_sc_hd__xnor2_1 _7174_ (.A(_2231_),
    .B(_2112_),
    .Y(_2232_));
 sky130_fd_sc_hd__xnor2_1 _7175_ (.A(_1191_),
    .B(_1193_),
    .Y(_2233_));
 sky130_fd_sc_hd__and2_1 _7176_ (.A(_1011_),
    .B(_1017_),
    .X(_2235_));
 sky130_fd_sc_hd__or2_1 _7177_ (.A(_1018_),
    .B(_2235_),
    .X(_2236_));
 sky130_fd_sc_hd__xnor2_1 _7178_ (.A(_2064_),
    .B(_2109_),
    .Y(_2237_));
 sky130_fd_sc_hd__nor2_1 _7179_ (.A(_2236_),
    .B(_2237_),
    .Y(_2238_));
 sky130_fd_sc_hd__a22o_1 _7180_ (.A1(_0726_),
    .A2(_4142_),
    .B1(_4210_),
    .B2(_0730_),
    .X(_2239_));
 sky130_fd_sc_hd__o21a_1 _7181_ (.A1(_1013_),
    .A2(_1015_),
    .B1(_2239_),
    .X(_2240_));
 sky130_fd_sc_hd__o21bai_1 _7182_ (.A1(_2080_),
    .A2(_2101_),
    .B1_N(_1015_),
    .Y(_2241_));
 sky130_fd_sc_hd__a21oi_1 _7183_ (.A1(_2080_),
    .A2(_2101_),
    .B1(_2241_),
    .Y(_2242_));
 sky130_fd_sc_hd__nand2_1 _7184_ (.A(_2076_),
    .B(_2103_),
    .Y(_2243_));
 sky130_fd_sc_hd__or2_1 _7185_ (.A(_2076_),
    .B(_2103_),
    .X(_2244_));
 sky130_fd_sc_hd__a22o_1 _7186_ (.A1(_2240_),
    .A2(_2242_),
    .B1(_2243_),
    .B2(_2244_),
    .X(_2245_));
 sky130_fd_sc_hd__o21ai_1 _7187_ (.A1(_2240_),
    .A2(_2242_),
    .B1(_2245_),
    .Y(_2246_));
 sky130_fd_sc_hd__xnor2_1 _7188_ (.A(_2070_),
    .B(_2105_),
    .Y(_2247_));
 sky130_fd_sc_hd__nand3_1 _7189_ (.A(_1000_),
    .B(_1014_),
    .C(_1016_),
    .Y(_2248_));
 sky130_fd_sc_hd__o2bb2a_1 _7190_ (.A1_N(_1017_),
    .A2_N(_2248_),
    .B1(_2247_),
    .B2(_2246_),
    .X(_2249_));
 sky130_fd_sc_hd__a221oi_1 _7191_ (.A1(_2236_),
    .A2(_2237_),
    .B1(_2246_),
    .B2(_2247_),
    .C1(_2249_),
    .Y(_2250_));
 sky130_fd_sc_hd__o22a_1 _7192_ (.A1(_2232_),
    .A2(_2233_),
    .B1(_2238_),
    .B2(_2250_),
    .X(_2251_));
 sky130_fd_sc_hd__xnor2_1 _7193_ (.A(_2052_),
    .B(_2114_),
    .Y(_2252_));
 sky130_fd_sc_hd__and2_1 _7194_ (.A(_1190_),
    .B(_1194_),
    .X(_2253_));
 sky130_fd_sc_hd__or2_1 _7195_ (.A(_1195_),
    .B(_2253_),
    .X(_2254_));
 sky130_fd_sc_hd__a2bb2o_1 _7196_ (.A1_N(_2252_),
    .A2_N(_2254_),
    .B1(_2232_),
    .B2(_2233_),
    .X(_2256_));
 sky130_fd_sc_hd__a22o_1 _7197_ (.A1(_2228_),
    .A2(_2229_),
    .B1(_2252_),
    .B2(_2254_),
    .X(_2257_));
 sky130_fd_sc_hd__o21bai_1 _7198_ (.A1(_2251_),
    .A2(_2256_),
    .B1_N(_2257_),
    .Y(_2258_));
 sky130_fd_sc_hd__and2_1 _7199_ (.A(_2224_),
    .B(_2226_),
    .X(_2259_));
 sky130_fd_sc_hd__a31oi_2 _7200_ (.A1(_2227_),
    .A2(_2230_),
    .A3(_2258_),
    .B1(_2259_),
    .Y(_2260_));
 sky130_fd_sc_hd__nor2_1 _7201_ (.A(_2220_),
    .B(_2222_),
    .Y(_2261_));
 sky130_fd_sc_hd__a21o_1 _7202_ (.A1(_2223_),
    .A2(_2260_),
    .B1(_2261_),
    .X(_2262_));
 sky130_fd_sc_hd__and3_1 _7203_ (.A(_1206_),
    .B(_2216_),
    .C(_2217_),
    .X(_2263_));
 sky130_fd_sc_hd__a21o_1 _7204_ (.A1(_2219_),
    .A2(_2262_),
    .B1(_2263_),
    .X(_2264_));
 sky130_fd_sc_hd__nor2_1 _7205_ (.A(_2211_),
    .B(_2214_),
    .Y(_2265_));
 sky130_fd_sc_hd__a21o_1 _7206_ (.A1(_2215_),
    .A2(_2264_),
    .B1(_2265_),
    .X(_2266_));
 sky130_fd_sc_hd__and2_1 _7207_ (.A(_2207_),
    .B(_2209_),
    .X(_2267_));
 sky130_fd_sc_hd__a21o_1 _7208_ (.A1(_2210_),
    .A2(_2266_),
    .B1(_2267_),
    .X(_2268_));
 sky130_fd_sc_hd__and2b_1 _7209_ (.A_N(_2202_),
    .B(_2204_),
    .X(_2269_));
 sky130_fd_sc_hd__a21o_1 _7210_ (.A1(_2205_),
    .A2(_2268_),
    .B1(_2269_),
    .X(_2270_));
 sky130_fd_sc_hd__nor2_1 _7211_ (.A(_2199_),
    .B(_2200_),
    .Y(_2271_));
 sky130_fd_sc_hd__a21o_1 _7212_ (.A1(_2201_),
    .A2(_2270_),
    .B1(_2271_),
    .X(_2272_));
 sky130_fd_sc_hd__nor2_1 _7213_ (.A(_2194_),
    .B(_2196_),
    .Y(_2273_));
 sky130_fd_sc_hd__a21oi_4 _7214_ (.A1(_2272_),
    .A2(_2197_),
    .B1(_2273_),
    .Y(_2274_));
 sky130_fd_sc_hd__or2_1 _7215_ (.A(_2188_),
    .B(_2191_),
    .X(_2275_));
 sky130_fd_sc_hd__o21ai_4 _7216_ (.A1(_2274_),
    .A2(_2193_),
    .B1(_2275_),
    .Y(_2277_));
 sky130_fd_sc_hd__and3_1 _7217_ (.A(_2002_),
    .B(_2007_),
    .C(_2147_),
    .X(_2278_));
 sky130_fd_sc_hd__a21oi_2 _7218_ (.A1(_2007_),
    .A2(_2147_),
    .B1(_2002_),
    .Y(_2279_));
 sky130_fd_sc_hd__nor2_4 _7219_ (.A(_2279_),
    .B(_2278_),
    .Y(_2280_));
 sky130_fd_sc_hd__a21oi_1 _7220_ (.A1(_1141_),
    .A2(_1219_),
    .B1(_1220_),
    .Y(_2281_));
 sky130_fd_sc_hd__and3_1 _7221_ (.A(_1220_),
    .B(_1141_),
    .C(_1219_),
    .X(_2282_));
 sky130_fd_sc_hd__nor2_1 _7222_ (.A(_2281_),
    .B(_2282_),
    .Y(_2283_));
 sky130_fd_sc_hd__xor2_2 _7223_ (.A(_2280_),
    .B(_2283_),
    .X(_2284_));
 sky130_fd_sc_hd__and2_1 _7224_ (.A(_2280_),
    .B(_2283_),
    .X(_2285_));
 sky130_fd_sc_hd__a21o_1 _7225_ (.A1(_2284_),
    .A2(_2277_),
    .B1(_2285_),
    .X(_2286_));
 sky130_fd_sc_hd__xnor2_2 _7226_ (.A(_1997_),
    .B(_2149_),
    .Y(_2288_));
 sky130_fd_sc_hd__and3_1 _7227_ (.A(_1222_),
    .B(_1136_),
    .C(_1221_),
    .X(_2289_));
 sky130_fd_sc_hd__or2_1 _7228_ (.A(_1223_),
    .B(_2289_),
    .X(_2290_));
 sky130_fd_sc_hd__nor2_1 _7229_ (.A(_2288_),
    .B(_2290_),
    .Y(_2291_));
 sky130_fd_sc_hd__and2_1 _7230_ (.A(_2288_),
    .B(_2290_),
    .X(_2292_));
 sky130_fd_sc_hd__nor2_1 _7231_ (.A(_2291_),
    .B(_2292_),
    .Y(_2293_));
 sky130_fd_sc_hd__a21o_1 _7232_ (.A1(_2293_),
    .A2(_2286_),
    .B1(_2291_),
    .X(_2294_));
 sky130_fd_sc_hd__and2b_1 _7233_ (.A_N(_2183_),
    .B(_2185_),
    .X(_2295_));
 sky130_fd_sc_hd__a21o_1 _7234_ (.A1(_2294_),
    .A2(_2186_),
    .B1(_2295_),
    .X(_2296_));
 sky130_fd_sc_hd__a21o_1 _7235_ (.A1(_2296_),
    .A2(_2182_),
    .B1(_2180_),
    .X(_2297_));
 sky130_fd_sc_hd__and2_1 _7236_ (.A(_2166_),
    .B(_2168_),
    .X(_2298_));
 sky130_fd_sc_hd__a211o_1 _7237_ (.A1(_2297_),
    .A2(_2176_),
    .B1(_2298_),
    .C1(_2174_),
    .X(_2299_));
 sky130_fd_sc_hd__and2_1 _7238_ (.A(_2157_),
    .B(_2158_),
    .X(_2300_));
 sky130_fd_sc_hd__and3_1 _7239_ (.A(_1233_),
    .B(_1113_),
    .C(_1232_),
    .X(_2301_));
 sky130_fd_sc_hd__or2_1 _7240_ (.A(_1234_),
    .B(_2301_),
    .X(_2302_));
 sky130_fd_sc_hd__o21a_1 _7241_ (.A1(_2159_),
    .A2(_2300_),
    .B1(_2302_),
    .X(_2303_));
 sky130_fd_sc_hd__nor3_1 _7242_ (.A(_2159_),
    .B(_2300_),
    .C(_2302_),
    .Y(_2304_));
 sky130_fd_sc_hd__nor2_2 _7243_ (.A(_2303_),
    .B(_2304_),
    .Y(_2305_));
 sky130_fd_sc_hd__a31o_1 _7244_ (.A1(_2305_),
    .A2(_2299_),
    .A3(_2169_),
    .B1(_2304_),
    .X(_2306_));
 sky130_fd_sc_hd__nand4_1 _7245_ (.A(_1345_),
    .B(_1611_),
    .C(_2160_),
    .D(_2163_),
    .Y(_2307_));
 sky130_fd_sc_hd__and3_1 _7246_ (.A(_1239_),
    .B(_1098_),
    .C(_1238_),
    .X(_2309_));
 sky130_fd_sc_hd__nor2_1 _7247_ (.A(_1240_),
    .B(_2309_),
    .Y(_2310_));
 sky130_fd_sc_hd__or3_1 _7248_ (.A(_1103_),
    .B(_1236_),
    .C(_1237_),
    .X(_2311_));
 sky130_fd_sc_hd__and2_1 _7249_ (.A(_1238_),
    .B(_2311_),
    .X(_2312_));
 sky130_fd_sc_hd__o2111ai_2 _7250_ (.A1(_2164_),
    .A2(_2306_),
    .B1(_2307_),
    .C1(_2310_),
    .D1(_2312_),
    .Y(_2313_));
 sky130_fd_sc_hd__nor3_1 _7251_ (.A(_1093_),
    .B(_1240_),
    .C(_1241_),
    .Y(_2314_));
 sky130_fd_sc_hd__or2_1 _7252_ (.A(_1242_),
    .B(_2314_),
    .X(_2315_));
 sky130_fd_sc_hd__xnor2_1 _7253_ (.A(_1085_),
    .B(_1243_),
    .Y(_2316_));
 sky130_fd_sc_hd__or3_4 _7254_ (.A(_2316_),
    .B(_2315_),
    .C(_2313_),
    .X(_2317_));
 sky130_fd_sc_hd__and2b_1 _7255_ (.A_N(_1246_),
    .B(_1245_),
    .X(_2318_));
 sky130_fd_sc_hd__or2_4 _7256_ (.A(_1247_),
    .B(_2318_),
    .X(_2319_));
 sky130_fd_sc_hd__xor2_1 _7257_ (.A(_1247_),
    .B(_1249_),
    .X(_2320_));
 sky130_fd_sc_hd__nor3b_4 _7258_ (.A(_2319_),
    .B(_2317_),
    .C_N(_2320_),
    .Y(_2321_));
 sky130_fd_sc_hd__or3_1 _7259_ (.A(_0550_),
    .B(_0716_),
    .C(_0717_),
    .X(_2322_));
 sky130_fd_sc_hd__and2_1 _7260_ (.A(_0718_),
    .B(_2322_),
    .X(_2323_));
 sky130_fd_sc_hd__o21ai_2 _7261_ (.A1(_2321_),
    .A2(_1250_),
    .B1(_2323_),
    .Y(_2324_));
 sky130_fd_sc_hd__nand2_1 _7262_ (.A(_0187_),
    .B(_0323_),
    .Y(_2325_));
 sky130_fd_sc_hd__or2b_1 _7263_ (.A(_2325_),
    .B_N(_0324_),
    .X(_2326_));
 sky130_fd_sc_hd__nand2_1 _7264_ (.A(_0325_),
    .B(_2326_),
    .Y(_2327_));
 sky130_fd_sc_hd__a31oi_2 _7265_ (.A1(_0456_),
    .A2(_0718_),
    .A3(_2324_),
    .B1(_2327_),
    .Y(_2328_));
 sky130_fd_sc_hd__and4_1 _7266_ (.A(_2324_),
    .B(_0456_),
    .C(_0718_),
    .D(_2327_),
    .X(_2330_));
 sky130_fd_sc_hd__or2_4 _7267_ (.A(_2328_),
    .B(_2330_),
    .X(_2331_));
 sky130_fd_sc_hd__nand3_1 _7268_ (.A(_0322_),
    .B(_0190_),
    .C(_0320_),
    .Y(_2332_));
 sky130_fd_sc_hd__and2_1 _7269_ (.A(_0323_),
    .B(_2332_),
    .X(_2333_));
 sky130_fd_sc_hd__or3_4 _7270_ (.A(_1250_),
    .B(_2321_),
    .C(_2323_),
    .X(_2334_));
 sky130_fd_sc_hd__and2_4 _7271_ (.A(_2334_),
    .B(_2324_),
    .X(_2335_));
 sky130_fd_sc_hd__xnor2_2 _7272_ (.A(_2333_),
    .B(_2335_),
    .Y(_2336_));
 sky130_fd_sc_hd__or2_4 _7273_ (.A(_2336_),
    .B(_2331_),
    .X(_2337_));
 sky130_fd_sc_hd__nor2_1 _7274_ (.A(_2317_),
    .B(_2319_),
    .Y(_2338_));
 sky130_fd_sc_hd__xor2_1 _7275_ (.A(_2338_),
    .B(_2320_),
    .X(_2339_));
 sky130_fd_sc_hd__or3_1 _7276_ (.A(_0319_),
    .B(_0195_),
    .C(_0317_),
    .X(_2340_));
 sky130_fd_sc_hd__and2_1 _7277_ (.A(_0320_),
    .B(_2340_),
    .X(_2341_));
 sky130_fd_sc_hd__nor2_1 _7278_ (.A(_2339_),
    .B(_2341_),
    .Y(_2342_));
 sky130_fd_sc_hd__nand2_2 _7279_ (.A(net105),
    .B(_2319_),
    .Y(_2343_));
 sky130_fd_sc_hd__nand2b_4 _7280_ (.A_N(_2338_),
    .B(_2343_),
    .Y(_2344_));
 sky130_fd_sc_hd__xnor2_2 _7281_ (.A(_0197_),
    .B(_0316_),
    .Y(_2345_));
 sky130_fd_sc_hd__and2b_1 _7282_ (.A_N(_2344_),
    .B(_2345_),
    .X(_2346_));
 sky130_fd_sc_hd__and2_1 _7283_ (.A(_2339_),
    .B(_2341_),
    .X(_2347_));
 sky130_fd_sc_hd__or2_1 _7284_ (.A(_2346_),
    .B(_2347_),
    .X(_2348_));
 sky130_fd_sc_hd__nor3b_2 _7285_ (.A(_2337_),
    .B(_2342_),
    .C_N(_2348_),
    .Y(_2349_));
 sky130_fd_sc_hd__or2_1 _7286_ (.A(_2313_),
    .B(_2315_),
    .X(_2351_));
 sky130_fd_sc_hd__nand2_1 _7287_ (.A(_2351_),
    .B(_2316_),
    .Y(_2352_));
 sky130_fd_sc_hd__nor3_1 _7288_ (.A(_0314_),
    .B(_0206_),
    .C(_0313_),
    .Y(_2353_));
 sky130_fd_sc_hd__nor2_1 _7289_ (.A(_0315_),
    .B(_2353_),
    .Y(_2354_));
 sky130_fd_sc_hd__a21oi_1 _7290_ (.A1(_2317_),
    .A2(_2352_),
    .B1(_2354_),
    .Y(_2355_));
 sky130_fd_sc_hd__and2_4 _7291_ (.A(_2307_),
    .B(_2306_),
    .X(_2356_));
 sky130_fd_sc_hd__o21a_1 _7292_ (.A1(_2164_),
    .A2(_2356_),
    .B1(_2312_),
    .X(_2357_));
 sky130_fd_sc_hd__xor2_1 _7293_ (.A(_2310_),
    .B(_2357_),
    .X(_2358_));
 sky130_fd_sc_hd__nor3_1 _7294_ (.A(_0309_),
    .B(_0216_),
    .C(_0307_),
    .Y(_2359_));
 sky130_fd_sc_hd__nor2_1 _7295_ (.A(_0310_),
    .B(_2359_),
    .Y(_2360_));
 sky130_fd_sc_hd__nor2_1 _7296_ (.A(_2358_),
    .B(_2360_),
    .Y(_2361_));
 sky130_fd_sc_hd__and3_1 _7297_ (.A(_0303_),
    .B(_0226_),
    .C(_0301_),
    .X(_2362_));
 sky130_fd_sc_hd__or2_1 _7298_ (.A(_0304_),
    .B(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__and2b_1 _7299_ (.A_N(_2164_),
    .B(_2307_),
    .X(_2364_));
 sky130_fd_sc_hd__xnor2_1 _7300_ (.A(_2306_),
    .B(_2364_),
    .Y(_2365_));
 sky130_fd_sc_hd__nor2_1 _7301_ (.A(_2363_),
    .B(_2365_),
    .Y(_2366_));
 sky130_fd_sc_hd__and2_1 _7302_ (.A(_2363_),
    .B(_2365_),
    .X(_2367_));
 sky130_fd_sc_hd__or2_4 _7303_ (.A(_2366_),
    .B(_2367_),
    .X(_2368_));
 sky130_fd_sc_hd__nand3_1 _7304_ (.A(_0300_),
    .B(_0231_),
    .C(_0298_),
    .Y(_2369_));
 sky130_fd_sc_hd__and2_1 _7305_ (.A(_0301_),
    .B(_2369_),
    .X(_2370_));
 sky130_fd_sc_hd__nand2_1 _7306_ (.A(_2169_),
    .B(_2299_),
    .Y(_2372_));
 sky130_fd_sc_hd__xnor2_1 _7307_ (.A(_2372_),
    .B(_2305_),
    .Y(_2373_));
 sky130_fd_sc_hd__xor2_1 _7308_ (.A(_2370_),
    .B(_2373_),
    .X(_2374_));
 sky130_fd_sc_hd__nand3_1 _7309_ (.A(_0297_),
    .B(_0236_),
    .C(_0295_),
    .Y(_2375_));
 sky130_fd_sc_hd__nand2_1 _7310_ (.A(_0298_),
    .B(_2375_),
    .Y(_2376_));
 sky130_fd_sc_hd__a21o_1 _7311_ (.A1(_2176_),
    .A2(_2297_),
    .B1(_2174_),
    .X(_2377_));
 sky130_fd_sc_hd__and2b_1 _7312_ (.A_N(_2298_),
    .B(_2169_),
    .X(_2378_));
 sky130_fd_sc_hd__xnor2_1 _7313_ (.A(_2377_),
    .B(_2378_),
    .Y(_2379_));
 sky130_fd_sc_hd__nand2_1 _7314_ (.A(_2376_),
    .B(_2379_),
    .Y(_2380_));
 sky130_fd_sc_hd__xor2_1 _7315_ (.A(_2176_),
    .B(_2297_),
    .X(_2381_));
 sky130_fd_sc_hd__or3_1 _7316_ (.A(_0294_),
    .B(_0240_),
    .C(_0292_),
    .X(_2382_));
 sky130_fd_sc_hd__and2_1 _7317_ (.A(_0295_),
    .B(_2382_),
    .X(_2383_));
 sky130_fd_sc_hd__xor2_1 _7318_ (.A(_2381_),
    .B(_2383_),
    .X(_2384_));
 sky130_fd_sc_hd__xnor2_2 _7319_ (.A(_2182_),
    .B(_2296_),
    .Y(_2385_));
 sky130_fd_sc_hd__nor3_1 _7320_ (.A(_0291_),
    .B(_0245_),
    .C(_0289_),
    .Y(_2386_));
 sky130_fd_sc_hd__nor2_1 _7321_ (.A(_0292_),
    .B(_2386_),
    .Y(_2387_));
 sky130_fd_sc_hd__xnor2_2 _7322_ (.A(_2385_),
    .B(_2387_),
    .Y(_2388_));
 sky130_fd_sc_hd__xnor2_2 _7323_ (.A(_2186_),
    .B(_2294_),
    .Y(_2389_));
 sky130_fd_sc_hd__and3_1 _7324_ (.A(_0288_),
    .B(_0248_),
    .C(_0286_),
    .X(_2390_));
 sky130_fd_sc_hd__or2_1 _7325_ (.A(_0289_),
    .B(_2390_),
    .X(_2391_));
 sky130_fd_sc_hd__xor2_2 _7326_ (.A(_2389_),
    .B(_2391_),
    .X(_2393_));
 sky130_fd_sc_hd__or3_1 _7327_ (.A(_0285_),
    .B(_0253_),
    .C(_0283_),
    .X(_2394_));
 sky130_fd_sc_hd__and2_1 _7328_ (.A(_0286_),
    .B(_2394_),
    .X(_2395_));
 sky130_fd_sc_hd__inv_2 _7329_ (.A(_2395_),
    .Y(_2396_));
 sky130_fd_sc_hd__xnor2_1 _7330_ (.A(_2286_),
    .B(_2293_),
    .Y(_2397_));
 sky130_fd_sc_hd__nand2_1 _7331_ (.A(_2396_),
    .B(_2397_),
    .Y(_2398_));
 sky130_fd_sc_hd__xnor2_2 _7332_ (.A(_2193_),
    .B(_2274_),
    .Y(_2399_));
 sky130_fd_sc_hd__or3_1 _7333_ (.A(_0263_),
    .B(_0277_),
    .C(_0278_),
    .X(_2400_));
 sky130_fd_sc_hd__and2_1 _7334_ (.A(_0279_),
    .B(_2400_),
    .X(_2401_));
 sky130_fd_sc_hd__xnor2_2 _7335_ (.A(_2399_),
    .B(_2401_),
    .Y(_2402_));
 sky130_fd_sc_hd__xnor2_1 _7336_ (.A(_2197_),
    .B(_2272_),
    .Y(_2404_));
 sky130_fd_sc_hd__xnor2_1 _7337_ (.A(_0274_),
    .B(_0276_),
    .Y(_2405_));
 sky130_fd_sc_hd__nand2_1 _7338_ (.A(_2404_),
    .B(_2405_),
    .Y(_2406_));
 sky130_fd_sc_hd__xor2_1 _7339_ (.A(_2201_),
    .B(_2270_),
    .X(_2407_));
 sky130_fd_sc_hd__xnor2_1 _7340_ (.A(_0266_),
    .B(_0271_),
    .Y(_2408_));
 sky130_fd_sc_hd__xor2_1 _7341_ (.A(_2205_),
    .B(_2268_),
    .X(_2409_));
 sky130_fd_sc_hd__a21oi_1 _7342_ (.A1(_4210_),
    .A2(_4111_),
    .B1(_0265_),
    .Y(_2410_));
 sky130_fd_sc_hd__nor2_1 _7343_ (.A(_0266_),
    .B(_2410_),
    .Y(_2411_));
 sky130_fd_sc_hd__xnor2_1 _7344_ (.A(_2210_),
    .B(_2266_),
    .Y(_2412_));
 sky130_fd_sc_hd__and2_1 _7345_ (.A(_4032_),
    .B(_4034_),
    .X(_2413_));
 sky130_fd_sc_hd__or2_1 _7346_ (.A(_4035_),
    .B(_2413_),
    .X(_2415_));
 sky130_fd_sc_hd__nor2_1 _7347_ (.A(_2412_),
    .B(_2415_),
    .Y(_2416_));
 sky130_fd_sc_hd__nand2_1 _7348_ (.A(_2219_),
    .B(_2262_),
    .Y(_2417_));
 sky130_fd_sc_hd__xor2_1 _7349_ (.A(_2223_),
    .B(_2260_),
    .X(_2418_));
 sky130_fd_sc_hd__a22oi_1 _7350_ (.A1(_4142_),
    .A2(_2546_),
    .B1(_2458_),
    .B2(_4210_),
    .Y(_2419_));
 sky130_fd_sc_hd__nor2_1 _7351_ (.A(_3566_),
    .B(_2419_),
    .Y(_2420_));
 sky130_fd_sc_hd__a31o_1 _7352_ (.A1(_4210_),
    .A2(_2546_),
    .A3(_2418_),
    .B1(_2420_),
    .X(_2421_));
 sky130_fd_sc_hd__or2_1 _7353_ (.A(_2219_),
    .B(_2262_),
    .X(_2422_));
 sky130_fd_sc_hd__and4_1 _7354_ (.A(_4210_),
    .B(_2546_),
    .C(_2420_),
    .D(_2418_),
    .X(_2423_));
 sky130_fd_sc_hd__a31o_1 _7355_ (.A1(_2417_),
    .A2(_2421_),
    .A3(_2422_),
    .B1(_2423_),
    .X(_2424_));
 sky130_fd_sc_hd__xnor2_1 _7356_ (.A(_3871_),
    .B(_4031_),
    .Y(_2426_));
 sky130_fd_sc_hd__or2_1 _7357_ (.A(_2215_),
    .B(_2264_),
    .X(_2427_));
 sky130_fd_sc_hd__nand2_1 _7358_ (.A(_2215_),
    .B(_2264_),
    .Y(_2428_));
 sky130_fd_sc_hd__a22o_1 _7359_ (.A1(_2424_),
    .A2(_2426_),
    .B1(_2427_),
    .B2(_2428_),
    .X(_2429_));
 sky130_fd_sc_hd__nand2_1 _7360_ (.A(_2412_),
    .B(_2415_),
    .Y(_2430_));
 sky130_fd_sc_hd__o211a_1 _7361_ (.A1(_2424_),
    .A2(_2426_),
    .B1(_2429_),
    .C1(_2430_),
    .X(_2431_));
 sky130_fd_sc_hd__o22a_1 _7362_ (.A1(_2409_),
    .A2(_2411_),
    .B1(_2416_),
    .B2(_2431_),
    .X(_2432_));
 sky130_fd_sc_hd__a221o_1 _7363_ (.A1(_2407_),
    .A2(_2408_),
    .B1(_2409_),
    .B2(_2411_),
    .C1(_2432_),
    .X(_2433_));
 sky130_fd_sc_hd__or2_1 _7364_ (.A(_2407_),
    .B(_2408_),
    .X(_2434_));
 sky130_fd_sc_hd__nor2_1 _7365_ (.A(_2404_),
    .B(_2405_),
    .Y(_2435_));
 sky130_fd_sc_hd__a31o_2 _7366_ (.A1(_2406_),
    .A2(_2433_),
    .A3(_2434_),
    .B1(_2435_),
    .X(_2437_));
 sky130_fd_sc_hd__and2b_1 _7367_ (.A_N(_2399_),
    .B(_2401_),
    .X(_2438_));
 sky130_fd_sc_hd__a21o_1 _7368_ (.A1(_2402_),
    .A2(_2437_),
    .B1(_2438_),
    .X(_2439_));
 sky130_fd_sc_hd__xnor2_2 _7369_ (.A(_2277_),
    .B(_2284_),
    .Y(_2440_));
 sky130_fd_sc_hd__or2_1 _7370_ (.A(_0280_),
    .B(_0282_),
    .X(_2441_));
 sky130_fd_sc_hd__and2b_1 _7371_ (.A_N(_0283_),
    .B(_2441_),
    .X(_2442_));
 sky130_fd_sc_hd__xnor2_2 _7372_ (.A(_2440_),
    .B(_2442_),
    .Y(_2443_));
 sky130_fd_sc_hd__and2b_1 _7373_ (.A_N(_2440_),
    .B(_2442_),
    .X(_2444_));
 sky130_fd_sc_hd__a21o_1 _7374_ (.A1(_2439_),
    .A2(_2443_),
    .B1(_2444_),
    .X(_2445_));
 sky130_fd_sc_hd__nor2_1 _7375_ (.A(_2396_),
    .B(_2397_),
    .Y(_2446_));
 sky130_fd_sc_hd__a21o_1 _7376_ (.A1(_2398_),
    .A2(_2445_),
    .B1(_2446_),
    .X(_2448_));
 sky130_fd_sc_hd__nor2_1 _7377_ (.A(_2389_),
    .B(_2391_),
    .Y(_2449_));
 sky130_fd_sc_hd__a21o_1 _7378_ (.A1(_2393_),
    .A2(_2448_),
    .B1(_2449_),
    .X(_2450_));
 sky130_fd_sc_hd__and2b_1 _7379_ (.A_N(_2385_),
    .B(_2387_),
    .X(_2451_));
 sky130_fd_sc_hd__a21o_1 _7380_ (.A1(_2388_),
    .A2(_2450_),
    .B1(_2451_),
    .X(_2452_));
 sky130_fd_sc_hd__and2_1 _7381_ (.A(_2381_),
    .B(_2383_),
    .X(_2453_));
 sky130_fd_sc_hd__a21o_1 _7382_ (.A1(_2384_),
    .A2(_2452_),
    .B1(_2453_),
    .X(_2454_));
 sky130_fd_sc_hd__nor2_1 _7383_ (.A(_2376_),
    .B(_2379_),
    .Y(_2455_));
 sky130_fd_sc_hd__a21o_1 _7384_ (.A1(_2380_),
    .A2(_2454_),
    .B1(_2455_),
    .X(_2456_));
 sky130_fd_sc_hd__and2_1 _7385_ (.A(_2370_),
    .B(_2373_),
    .X(_2457_));
 sky130_fd_sc_hd__a21oi_1 _7386_ (.A1(_2374_),
    .A2(_2456_),
    .B1(_2457_),
    .Y(_2459_));
 sky130_fd_sc_hd__o21bai_4 _7387_ (.A1(_2459_),
    .A2(_2368_),
    .B1_N(_2366_),
    .Y(_2460_));
 sky130_fd_sc_hd__nor3_1 _7388_ (.A(_2312_),
    .B(_2164_),
    .C(_2356_),
    .Y(_2461_));
 sky130_fd_sc_hd__or2_4 _7389_ (.A(_2461_),
    .B(_2357_),
    .X(_2462_));
 sky130_fd_sc_hd__or3b_1 _7390_ (.A(_0221_),
    .B(_0304_),
    .C_N(_0306_),
    .X(_2463_));
 sky130_fd_sc_hd__or2b_1 _7391_ (.A(_0307_),
    .B_N(_2463_),
    .X(_2464_));
 sky130_fd_sc_hd__xor2_2 _7392_ (.A(_2464_),
    .B(_2462_),
    .X(_2465_));
 sky130_fd_sc_hd__nor2_1 _7393_ (.A(_2462_),
    .B(_2464_),
    .Y(_2466_));
 sky130_fd_sc_hd__a21oi_2 _7394_ (.A1(_2465_),
    .A2(_2460_),
    .B1(_2466_),
    .Y(_2467_));
 sky130_fd_sc_hd__and2_1 _7395_ (.A(_2358_),
    .B(_2360_),
    .X(_2468_));
 sky130_fd_sc_hd__o21ba_4 _7396_ (.A1(_2361_),
    .A2(_2467_),
    .B1_N(_2468_),
    .X(_2470_));
 sky130_fd_sc_hd__nand2_1 _7397_ (.A(_2313_),
    .B(_2315_),
    .Y(_2471_));
 sky130_fd_sc_hd__nand2_1 _7398_ (.A(_2351_),
    .B(_2471_),
    .Y(_2472_));
 sky130_fd_sc_hd__nor3_1 _7399_ (.A(_0312_),
    .B(_0211_),
    .C(_0310_),
    .Y(_2473_));
 sky130_fd_sc_hd__nor2_1 _7400_ (.A(_0313_),
    .B(_2473_),
    .Y(_2474_));
 sky130_fd_sc_hd__xor2_2 _7401_ (.A(_2472_),
    .B(_2474_),
    .X(_2475_));
 sky130_fd_sc_hd__and3_1 _7402_ (.A(_2317_),
    .B(_2352_),
    .C(_2354_),
    .X(_2476_));
 sky130_fd_sc_hd__inv_2 _7403_ (.A(_2476_),
    .Y(_2477_));
 sky130_fd_sc_hd__or3_1 _7404_ (.A(_0313_),
    .B(_2472_),
    .C(_2473_),
    .X(_2478_));
 sky130_fd_sc_hd__o211a_4 _7405_ (.A1(_2475_),
    .A2(_2470_),
    .B1(_2477_),
    .C1(_2478_),
    .X(_2479_));
 sky130_fd_sc_hd__xnor2_2 _7406_ (.A(_2345_),
    .B(_2344_),
    .Y(_2481_));
 sky130_fd_sc_hd__nor2_1 _7407_ (.A(_2347_),
    .B(_2342_),
    .Y(_2482_));
 sky130_fd_sc_hd__nand2_1 _7408_ (.A(_2481_),
    .B(_2482_),
    .Y(_2483_));
 sky130_fd_sc_hd__nand2_1 _7409_ (.A(_2333_),
    .B(_2335_),
    .Y(_2484_));
 sky130_fd_sc_hd__or2_1 _7410_ (.A(_2330_),
    .B(_2484_),
    .X(_2485_));
 sky130_fd_sc_hd__o41ai_4 _7411_ (.A1(_2355_),
    .A2(_2479_),
    .A3(_2483_),
    .A4(_2337_),
    .B1(_2485_),
    .Y(_2486_));
 sky130_fd_sc_hd__xnor2_1 _7412_ (.A(_0326_),
    .B(_0179_),
    .Y(_2487_));
 sky130_fd_sc_hd__nand2_1 _7413_ (.A(_0177_),
    .B(_0327_),
    .Y(_2488_));
 sky130_fd_sc_hd__xnor2_1 _7414_ (.A(_2488_),
    .B(_0329_),
    .Y(_2489_));
 sky130_fd_sc_hd__o311a_4 _7415_ (.A1(_2328_),
    .A2(_2486_),
    .A3(_2349_),
    .B1(_2487_),
    .C1(_2489_),
    .X(_2490_));
 sky130_fd_sc_hd__a21o_1 _7416_ (.A1(_0173_),
    .A2(_0330_),
    .B1(_0357_),
    .X(_2492_));
 sky130_fd_sc_hd__nand2_1 _7417_ (.A(_0332_),
    .B(_0334_),
    .Y(_2493_));
 sky130_fd_sc_hd__or2_1 _7418_ (.A(_0349_),
    .B(_0352_),
    .X(_2494_));
 sky130_fd_sc_hd__o21bai_1 _7419_ (.A1(_0344_),
    .A2(_0346_),
    .B1_N(_0345_),
    .Y(_2495_));
 sky130_fd_sc_hd__and2_1 _7420_ (.A(_3907_),
    .B(_4245_),
    .X(_2496_));
 sky130_fd_sc_hd__nand2_1 _7421_ (.A(_3804_),
    .B(_2496_),
    .Y(_2497_));
 sky130_fd_sc_hd__or2_1 _7422_ (.A(_3804_),
    .B(_2496_),
    .X(_2498_));
 sky130_fd_sc_hd__nand2_1 _7423_ (.A(_2497_),
    .B(_2498_),
    .Y(_2499_));
 sky130_fd_sc_hd__xnor2_1 _7424_ (.A(_2495_),
    .B(_2499_),
    .Y(_2500_));
 sky130_fd_sc_hd__and3_1 _7425_ (.A(_4092_),
    .B(_4107_),
    .C(_4111_),
    .X(_2501_));
 sky130_fd_sc_hd__a21oi_1 _7426_ (.A1(_4092_),
    .A2(_4107_),
    .B1(_4111_),
    .Y(_2503_));
 sky130_fd_sc_hd__or2_1 _7427_ (.A(_2501_),
    .B(_2503_),
    .X(_2504_));
 sky130_fd_sc_hd__nand2_1 _7428_ (.A(_0339_),
    .B(_2504_),
    .Y(_2505_));
 sky130_fd_sc_hd__mux2_1 _7429_ (.A0(_2505_),
    .A1(_2504_),
    .S(_0341_),
    .X(_2506_));
 sky130_fd_sc_hd__xnor2_1 _7430_ (.A(_2500_),
    .B(_2506_),
    .Y(_2507_));
 sky130_fd_sc_hd__xnor2_1 _7431_ (.A(_2494_),
    .B(_2507_),
    .Y(_2508_));
 sky130_fd_sc_hd__xnor2_1 _7432_ (.A(_2493_),
    .B(_2508_),
    .Y(_2509_));
 sky130_fd_sc_hd__a21oi_1 _7433_ (.A1(_0355_),
    .A2(_2492_),
    .B1(_2509_),
    .Y(_2510_));
 sky130_fd_sc_hd__and3_1 _7434_ (.A(_0355_),
    .B(_2492_),
    .C(_2509_),
    .X(_2511_));
 sky130_fd_sc_hd__nor2_1 _7435_ (.A(_2510_),
    .B(_2511_),
    .Y(_2512_));
 sky130_fd_sc_hd__and2b_1 _7436_ (.A_N(_2507_),
    .B(_2494_),
    .X(_2514_));
 sky130_fd_sc_hd__a21oi_1 _7437_ (.A1(_2500_),
    .A2(_2506_),
    .B1(_2514_),
    .Y(_2515_));
 sky130_fd_sc_hd__nor2_1 _7438_ (.A(_0341_),
    .B(_2501_),
    .Y(_2516_));
 sky130_fd_sc_hd__and3_1 _7439_ (.A(_2497_),
    .B(_2495_),
    .C(_2498_),
    .X(_2517_));
 sky130_fd_sc_hd__inv_2 _7440_ (.A(_2517_),
    .Y(_2518_));
 sky130_fd_sc_hd__and3_1 _7441_ (.A(_4092_),
    .B(_3907_),
    .C(_4245_),
    .X(_2519_));
 sky130_fd_sc_hd__a21oi_1 _7442_ (.A1(_4092_),
    .A2(_4245_),
    .B1(_3907_),
    .Y(_2520_));
 sky130_fd_sc_hd__a211o_1 _7443_ (.A1(_2497_),
    .A2(_2518_),
    .B1(_2519_),
    .C1(_2520_),
    .X(_2521_));
 sky130_fd_sc_hd__o211ai_1 _7444_ (.A1(_2519_),
    .A2(_2520_),
    .B1(_2497_),
    .C1(_2518_),
    .Y(_2522_));
 sky130_fd_sc_hd__and2_1 _7445_ (.A(_2521_),
    .B(_2522_),
    .X(_2523_));
 sky130_fd_sc_hd__and3_1 _7446_ (.A(_4107_),
    .B(_2516_),
    .C(_2523_),
    .X(_2525_));
 sky130_fd_sc_hd__a21oi_1 _7447_ (.A1(_4107_),
    .A2(_2516_),
    .B1(_2523_),
    .Y(_2526_));
 sky130_fd_sc_hd__or2_1 _7448_ (.A(_2525_),
    .B(_2526_),
    .X(_2527_));
 sky130_fd_sc_hd__xnor2_1 _7449_ (.A(_2515_),
    .B(_2527_),
    .Y(_2528_));
 sky130_fd_sc_hd__a21oi_1 _7450_ (.A1(_2493_),
    .A2(_2508_),
    .B1(_2510_),
    .Y(_2529_));
 sky130_fd_sc_hd__or2_1 _7451_ (.A(_2528_),
    .B(_2529_),
    .X(_2530_));
 sky130_fd_sc_hd__nand2_1 _7452_ (.A(_2528_),
    .B(_2529_),
    .Y(_2531_));
 sky130_fd_sc_hd__and2_1 _7453_ (.A(_2530_),
    .B(_2531_),
    .X(_2532_));
 sky130_fd_sc_hd__and4_1 _7454_ (.A(_2490_),
    .B(_0358_),
    .C(_2512_),
    .D(_2532_),
    .X(_2533_));
 sky130_fd_sc_hd__nor2_1 _7455_ (.A(_2515_),
    .B(_2527_),
    .Y(_2534_));
 sky130_fd_sc_hd__nand2_1 _7456_ (.A(_4092_),
    .B(_4245_),
    .Y(_2536_));
 sky130_fd_sc_hd__or2_1 _7457_ (.A(_4092_),
    .B(_4245_),
    .X(_2537_));
 sky130_fd_sc_hd__nand2_1 _7458_ (.A(_2536_),
    .B(_2537_),
    .Y(_2538_));
 sky130_fd_sc_hd__a21o_1 _7459_ (.A1(_2536_),
    .A2(_2537_),
    .B1(_2496_),
    .X(_2539_));
 sky130_fd_sc_hd__mux2_1 _7460_ (.A0(_2538_),
    .A1(_2539_),
    .S(_2521_),
    .X(_2540_));
 sky130_fd_sc_hd__and2b_1 _7461_ (.A_N(_2516_),
    .B(_2540_),
    .X(_2541_));
 sky130_fd_sc_hd__and2b_1 _7462_ (.A_N(_2540_),
    .B(_2516_),
    .X(_2542_));
 sky130_fd_sc_hd__nor2_1 _7463_ (.A(_2541_),
    .B(_2542_),
    .Y(_2543_));
 sky130_fd_sc_hd__o21a_1 _7464_ (.A1(_2525_),
    .A2(_2534_),
    .B1(_2543_),
    .X(_2544_));
 sky130_fd_sc_hd__nor3_1 _7465_ (.A(_2543_),
    .B(_2525_),
    .C(_2534_),
    .Y(_2545_));
 sky130_fd_sc_hd__nor2_1 _7466_ (.A(_2544_),
    .B(_2545_),
    .Y(_2547_));
 sky130_fd_sc_hd__xnor2_2 _7467_ (.A(_2530_),
    .B(_2547_),
    .Y(_2548_));
 sky130_fd_sc_hd__o21ai_1 _7468_ (.A1(_2521_),
    .A2(_2538_),
    .B1(_2536_),
    .Y(_2549_));
 sky130_fd_sc_hd__and2b_1 _7469_ (.A_N(_2530_),
    .B(_2547_),
    .X(_2550_));
 sky130_fd_sc_hd__nor2_1 _7470_ (.A(_2541_),
    .B(_2544_),
    .Y(_2551_));
 sky130_fd_sc_hd__or3b_1 _7471_ (.A(_2549_),
    .B(_2550_),
    .C_N(_2551_),
    .X(_2552_));
 sky130_fd_sc_hd__a21o_4 _7472_ (.A1(_2548_),
    .A2(_2533_),
    .B1(_2552_),
    .X(_2553_));
 sky130_fd_sc_hd__or2_1 _7473_ (.A(\M1.ua1.fa1.b ),
    .B(\M1.ua1.fa1.a ),
    .X(_2554_));
 sky130_fd_sc_hd__nand2_1 _7474_ (.A(\M1.ua1.fa1.b ),
    .B(\M1.ua1.fa1.a ),
    .Y(_2555_));
 sky130_fd_sc_hd__nand2_1 _7475_ (.A(_2554_),
    .B(_2555_),
    .Y(_2556_));
 sky130_fd_sc_hd__xor2_2 _7476_ (.A(_2403_),
    .B(_2556_),
    .X(_2558_));
 sky130_fd_sc_hd__or2_1 _7477_ (.A(\M1.ua1.fa2.b ),
    .B(\M1.ua1.fa2.a ),
    .X(_2559_));
 sky130_fd_sc_hd__nand2_1 _7478_ (.A(\M1.ua1.fa2.b ),
    .B(\M1.ua1.fa2.a ),
    .Y(_2560_));
 sky130_fd_sc_hd__nand2_2 _7479_ (.A(_2559_),
    .B(_2560_),
    .Y(_2561_));
 sky130_fd_sc_hd__nor2_1 _7480_ (.A(\M1.ua1.fa1.b ),
    .B(\M1.ua1.fa1.a ),
    .Y(_2562_));
 sky130_fd_sc_hd__o21a_2 _7481_ (.A1(_2403_),
    .A2(_2562_),
    .B1(_2555_),
    .X(_2563_));
 sky130_fd_sc_hd__xor2_4 _7482_ (.A(_2561_),
    .B(_2563_),
    .X(_2564_));
 sky130_fd_sc_hd__or2_2 _7483_ (.A(\M1.ua1.fa3.b ),
    .B(\M1.ua1.fa3.a ),
    .X(_2565_));
 sky130_fd_sc_hd__nand2_1 _7484_ (.A(\M1.ua1.fa3.b ),
    .B(\M1.ua1.fa3.a ),
    .Y(_2566_));
 sky130_fd_sc_hd__nand2_1 _7485_ (.A(_2565_),
    .B(_2566_),
    .Y(_2567_));
 sky130_fd_sc_hd__nand2_1 _7486_ (.A(_2560_),
    .B(_2563_),
    .Y(_2569_));
 sky130_fd_sc_hd__and2_2 _7487_ (.A(_2559_),
    .B(_2569_),
    .X(_2570_));
 sky130_fd_sc_hd__xnor2_2 _7488_ (.A(_2567_),
    .B(_2570_),
    .Y(_2571_));
 sky130_fd_sc_hd__o2111a_4 _7489_ (.A1(_2414_),
    .A2(net128),
    .B1(_2558_),
    .C1(_2564_),
    .D1(_2571_),
    .X(_2572_));
 sky130_fd_sc_hd__or2_1 _7490_ (.A(\M1.ua1.fa4.b ),
    .B(\M1.ua1.fa4.a ),
    .X(_2573_));
 sky130_fd_sc_hd__nand2_1 _7491_ (.A(\M1.ua1.fa4.b ),
    .B(\M1.ua1.fa4.a ),
    .Y(_2574_));
 sky130_fd_sc_hd__nand2_2 _7492_ (.A(_2573_),
    .B(_2574_),
    .Y(_2575_));
 sky130_fd_sc_hd__a21boi_4 _7493_ (.A1(_2565_),
    .A2(_2570_),
    .B1_N(_2566_),
    .Y(_2576_));
 sky130_fd_sc_hd__xor2_4 _7494_ (.A(_2575_),
    .B(_2576_),
    .X(_2577_));
 sky130_fd_sc_hd__or2_1 _7495_ (.A(\M1.ua1.fa5.b ),
    .B(\M1.ua1.fa5.a ),
    .X(_2578_));
 sky130_fd_sc_hd__nand2_1 _7496_ (.A(\M1.ua1.fa5.b ),
    .B(\M1.ua1.fa5.a ),
    .Y(_2580_));
 sky130_fd_sc_hd__nand2_1 _7497_ (.A(_2578_),
    .B(_2580_),
    .Y(_2581_));
 sky130_fd_sc_hd__nand2_1 _7498_ (.A(_2574_),
    .B(_2576_),
    .Y(_2582_));
 sky130_fd_sc_hd__and2_1 _7499_ (.A(_2573_),
    .B(_2582_),
    .X(_2583_));
 sky130_fd_sc_hd__xnor2_1 _7500_ (.A(_2581_),
    .B(_2583_),
    .Y(_2584_));
 sky130_fd_sc_hd__nand3_4 _7501_ (.A(_2572_),
    .B(_2577_),
    .C(_2584_),
    .Y(_2585_));
 sky130_fd_sc_hd__or2_1 _7502_ (.A(\M1.ua1.fa6.b ),
    .B(\M1.ua1.fa6.a ),
    .X(_2586_));
 sky130_fd_sc_hd__nand2_1 _7503_ (.A(\M1.ua1.fa6.b ),
    .B(\M1.ua1.fa6.a ),
    .Y(_2587_));
 sky130_fd_sc_hd__nand2_1 _7504_ (.A(_2586_),
    .B(_2587_),
    .Y(_2588_));
 sky130_fd_sc_hd__a21boi_1 _7505_ (.A1(_2578_),
    .A2(_2583_),
    .B1_N(_2580_),
    .Y(_2589_));
 sky130_fd_sc_hd__xnor2_1 _7506_ (.A(_2588_),
    .B(_2589_),
    .Y(_2591_));
 sky130_fd_sc_hd__xnor2_4 _7507_ (.A(_2591_),
    .B(_2585_),
    .Y(_2592_));
 sky130_fd_sc_hd__or2_4 _7508_ (.A(net87),
    .B(_2592_),
    .X(_2593_));
 sky130_fd_sc_hd__nand2_1 _7509_ (.A(net87),
    .B(_2592_),
    .Y(_2594_));
 sky130_fd_sc_hd__and2_1 _7510_ (.A(_2593_),
    .B(_2594_),
    .X(_2595_));
 sky130_fd_sc_hd__buf_6 _7511_ (.A(_2595_),
    .X(_2596_));
 sky130_fd_sc_hd__a21o_1 _7512_ (.A1(_2572_),
    .A2(_2577_),
    .B1(_2584_),
    .X(_2597_));
 sky130_fd_sc_hd__a21boi_2 _7513_ (.A1(_2585_),
    .A2(_2597_),
    .B1_N(net86),
    .Y(_2598_));
 sky130_fd_sc_hd__and3b_2 _7514_ (.A_N(net86),
    .B(_2585_),
    .C(_2597_),
    .X(_2599_));
 sky130_fd_sc_hd__xnor2_4 _7515_ (.A(_2572_),
    .B(_2577_),
    .Y(_2600_));
 sky130_fd_sc_hd__xor2_4 _7516_ (.A(net85),
    .B(_2600_),
    .X(_2602_));
 sky130_fd_sc_hd__nor3b_4 _7517_ (.A(_2598_),
    .B(_2599_),
    .C_N(_2602_),
    .Y(_2603_));
 sky130_fd_sc_hd__or3_1 _7518_ (.A(\M1.ua1.fa7.b ),
    .B(\M1.ua1.fa7.a ),
    .C(_2586_),
    .X(_2604_));
 sky130_fd_sc_hd__or3_1 _7519_ (.A(_2573_),
    .B(_2578_),
    .C(_2604_),
    .X(_2605_));
 sky130_fd_sc_hd__or3_1 _7520_ (.A(_2392_),
    .B(_2554_),
    .C(_2605_),
    .X(_2606_));
 sky130_fd_sc_hd__nor3_2 _7521_ (.A(_2559_),
    .B(_2565_),
    .C(_2606_),
    .Y(_2607_));
 sky130_fd_sc_hd__inv_2 _7522_ (.A(_2591_),
    .Y(_2608_));
 sky130_fd_sc_hd__and4_1 _7523_ (.A(_2572_),
    .B(_2577_),
    .C(_2584_),
    .D(_2608_),
    .X(_2609_));
 sky130_fd_sc_hd__xor2_1 _7524_ (.A(\M1.ua1.fa7.b ),
    .B(\M1.ua1.fa7.a ),
    .X(_2610_));
 sky130_fd_sc_hd__nand2_1 _7525_ (.A(_2587_),
    .B(_2589_),
    .Y(_2611_));
 sky130_fd_sc_hd__and2_1 _7526_ (.A(_2586_),
    .B(_2611_),
    .X(_2613_));
 sky130_fd_sc_hd__xnor2_1 _7527_ (.A(_2610_),
    .B(_2613_),
    .Y(_2614_));
 sky130_fd_sc_hd__xnor2_2 _7528_ (.A(_2614_),
    .B(_2609_),
    .Y(_2615_));
 sky130_fd_sc_hd__o21ai_4 _7529_ (.A1(_2607_),
    .A2(net114),
    .B1(net89),
    .Y(_2616_));
 sky130_fd_sc_hd__or3_4 _7530_ (.A(net89),
    .B(_2607_),
    .C(_2615_),
    .X(_2617_));
 sky130_fd_sc_hd__and2_4 _7531_ (.A(_2616_),
    .B(_2617_),
    .X(_2618_));
 sky130_fd_sc_hd__buf_8 _7532_ (.A(_2553_),
    .X(_2619_));
 sky130_fd_sc_hd__o211a_1 _7533_ (.A1(_2414_),
    .A2(_2619_),
    .B1(_2558_),
    .C1(_2564_),
    .X(_2620_));
 sky130_fd_sc_hd__xnor2_2 _7534_ (.A(_2620_),
    .B(_2571_),
    .Y(_2621_));
 sky130_fd_sc_hd__nor2_1 _7535_ (.A(net84),
    .B(_2621_),
    .Y(_2622_));
 sky130_fd_sc_hd__nand2_1 _7536_ (.A(net84),
    .B(_2621_),
    .Y(_2624_));
 sky130_fd_sc_hd__nand2b_4 _7537_ (.A_N(_2622_),
    .B(_2624_),
    .Y(_2625_));
 sky130_fd_sc_hd__inv_2 _7538_ (.A(net83),
    .Y(_2626_));
 sky130_fd_sc_hd__o21ai_4 _7539_ (.A1(_2619_),
    .A2(_2414_),
    .B1(_2558_),
    .Y(_2627_));
 sky130_fd_sc_hd__xnor2_4 _7540_ (.A(_2564_),
    .B(_2627_),
    .Y(_2628_));
 sky130_fd_sc_hd__xnor2_4 _7541_ (.A(_2626_),
    .B(_2628_),
    .Y(_2629_));
 sky130_fd_sc_hd__or3_1 _7542_ (.A(_2559_),
    .B(_2565_),
    .C(_2606_),
    .X(_2630_));
 sky130_fd_sc_hd__xnor2_1 _7543_ (.A(_2414_),
    .B(_2619_),
    .Y(_2631_));
 sky130_fd_sc_hd__and2_2 _7544_ (.A(_2630_),
    .B(_2631_),
    .X(_2632_));
 sky130_fd_sc_hd__xnor2_4 _7545_ (.A(net81),
    .B(_2632_),
    .Y(_2633_));
 sky130_fd_sc_hd__inv_2 _7546_ (.A(net82),
    .Y(_2635_));
 sky130_fd_sc_hd__o31a_1 _7547_ (.A1(_2414_),
    .A2(_2553_),
    .A3(_2558_),
    .B1(_2630_),
    .X(_2636_));
 sky130_fd_sc_hd__and3_1 _7548_ (.A(_2627_),
    .B(_2635_),
    .C(_2636_),
    .X(_2637_));
 sky130_fd_sc_hd__a21o_1 _7549_ (.A1(_2627_),
    .A2(_2636_),
    .B1(_2635_),
    .X(_2638_));
 sky130_fd_sc_hd__and2b_2 _7550_ (.A_N(net127),
    .B(_2638_),
    .X(_2639_));
 sky130_fd_sc_hd__and4bb_1 _7551_ (.A_N(_2625_),
    .B_N(_2629_),
    .C(_2639_),
    .D(_2633_),
    .X(_2640_));
 sky130_fd_sc_hd__and4_1 _7552_ (.A(_2618_),
    .B(_2603_),
    .C(_2596_),
    .D(_2640_),
    .X(_2641_));
 sky130_fd_sc_hd__buf_6 _7553_ (.A(_2641_),
    .X(_2642_));
 sky130_fd_sc_hd__nor2_1 _7554_ (.A(net85),
    .B(_2600_),
    .Y(_2643_));
 sky130_fd_sc_hd__nor2_1 _7555_ (.A(_2643_),
    .B(_2599_),
    .Y(_2644_));
 sky130_fd_sc_hd__xor2_1 _7556_ (.A(_2627_),
    .B(_2564_),
    .X(_2646_));
 sky130_fd_sc_hd__nor2_1 _7557_ (.A(net83),
    .B(_2646_),
    .Y(_2647_));
 sky130_fd_sc_hd__inv_2 _7558_ (.A(net81),
    .Y(_2648_));
 sky130_fd_sc_hd__a21o_1 _7559_ (.A1(_2630_),
    .A2(_2631_),
    .B1(_2648_),
    .X(_2649_));
 sky130_fd_sc_hd__o221a_1 _7560_ (.A1(_2626_),
    .A2(_2628_),
    .B1(_2649_),
    .B2(_2637_),
    .C1(_2638_),
    .X(_2650_));
 sky130_fd_sc_hd__o31a_1 _7561_ (.A1(_2622_),
    .A2(_2650_),
    .A3(_2647_),
    .B1(_2624_),
    .X(_2651_));
 sky130_fd_sc_hd__a2bb2o_4 _7562_ (.A1_N(_2598_),
    .A2_N(_2644_),
    .B1(_2603_),
    .B2(_2651_),
    .X(_2652_));
 sky130_fd_sc_hd__nand2_1 _7563_ (.A(_2593_),
    .B(_2617_),
    .Y(_2653_));
 sky130_fd_sc_hd__a21o_2 _7564_ (.A1(_2596_),
    .A2(_2652_),
    .B1(_2653_),
    .X(_2654_));
 sky130_fd_sc_hd__nand2_4 _7565_ (.A(_2616_),
    .B(_2654_),
    .Y(_2655_));
 sky130_fd_sc_hd__clkbuf_4 _7566_ (.A(_2655_),
    .X(_2657_));
 sky130_fd_sc_hd__buf_2 _7567_ (.A(_2657_),
    .X(_2658_));
 sky130_fd_sc_hd__o21a_2 _7568_ (.A1(_2607_),
    .A2(net114),
    .B1(net89),
    .X(_2659_));
 sky130_fd_sc_hd__a21oi_4 _7569_ (.A1(_2596_),
    .A2(_2652_),
    .B1(_2653_),
    .Y(_2660_));
 sky130_fd_sc_hd__nor2_2 _7570_ (.A(_2659_),
    .B(_2660_),
    .Y(_2661_));
 sky130_fd_sc_hd__or3_4 _7571_ (.A(_2659_),
    .B(_2660_),
    .C(_2641_),
    .X(_2662_));
 sky130_fd_sc_hd__buf_8 _7572_ (.A(_2662_),
    .X(_2663_));
 sky130_fd_sc_hd__a31o_1 _7573_ (.A1(_2648_),
    .A2(_2638_),
    .A3(_2632_),
    .B1(_2637_),
    .X(_2664_));
 sky130_fd_sc_hd__o211ai_1 _7574_ (.A1(net84),
    .A2(_2621_),
    .B1(_2646_),
    .C1(net83),
    .Y(_2665_));
 sky130_fd_sc_hd__o311a_1 _7575_ (.A1(_2622_),
    .A2(_2629_),
    .A3(_2664_),
    .B1(_2665_),
    .C1(_2624_),
    .X(_2666_));
 sky130_fd_sc_hd__or4_1 _7576_ (.A(_2659_),
    .B(_2651_),
    .C(_2660_),
    .D(_2642_),
    .X(_2668_));
 sky130_fd_sc_hd__a21bo_2 _7577_ (.A1(net131),
    .A2(_2666_),
    .B1_N(_2668_),
    .X(_2669_));
 sky130_fd_sc_hd__xor2_4 _7578_ (.A(net101),
    .B(_2669_),
    .X(_2670_));
 sky130_fd_sc_hd__nor2_2 _7579_ (.A(_2598_),
    .B(_2599_),
    .Y(_2671_));
 sky130_fd_sc_hd__nand2_1 _7580_ (.A(net85),
    .B(_2600_),
    .Y(_2672_));
 sky130_fd_sc_hd__a21o_1 _7581_ (.A1(_2672_),
    .A2(_2651_),
    .B1(_2643_),
    .X(_2673_));
 sky130_fd_sc_hd__o21ai_1 _7582_ (.A1(_2643_),
    .A2(_2666_),
    .B1(_2672_),
    .Y(_2674_));
 sky130_fd_sc_hd__mux2_2 _7583_ (.A0(_2673_),
    .A1(_2674_),
    .S(net131),
    .X(_2675_));
 sky130_fd_sc_hd__xnor2_4 _7584_ (.A(_2671_),
    .B(_2675_),
    .Y(_2676_));
 sky130_fd_sc_hd__and3_1 _7585_ (.A(_2661_),
    .B(_2670_),
    .C(_2676_),
    .X(_2677_));
 sky130_fd_sc_hd__buf_2 _7586_ (.A(_2677_),
    .X(_2679_));
 sky130_fd_sc_hd__buf_2 _7587_ (.A(_2679_),
    .X(_2680_));
 sky130_fd_sc_hd__nor2_1 _7588_ (.A(_2647_),
    .B(_2650_),
    .Y(_2681_));
 sky130_fd_sc_hd__nand2_1 _7589_ (.A(net83),
    .B(_2646_),
    .Y(_2682_));
 sky130_fd_sc_hd__o21a_1 _7590_ (.A1(_2647_),
    .A2(_2664_),
    .B1(_2682_),
    .X(_2683_));
 sky130_fd_sc_hd__mux2_4 _7591_ (.A0(_2681_),
    .A1(_2683_),
    .S(_2663_),
    .X(_2684_));
 sky130_fd_sc_hd__xor2_4 _7592_ (.A(_2625_),
    .B(_2684_),
    .X(_2685_));
 sky130_fd_sc_hd__clkbuf_4 _7593_ (.A(_2685_),
    .X(_2686_));
 sky130_fd_sc_hd__clkbuf_4 _7594_ (.A(_2686_),
    .X(_2687_));
 sky130_fd_sc_hd__o21ai_1 _7595_ (.A1(_2637_),
    .A2(_2649_),
    .B1(_2638_),
    .Y(_2688_));
 sky130_fd_sc_hd__mux2_4 _7596_ (.A0(_2688_),
    .A1(_2664_),
    .S(_2663_),
    .X(_2690_));
 sky130_fd_sc_hd__xnor2_4 _7597_ (.A(_2690_),
    .B(_2629_),
    .Y(_2691_));
 sky130_fd_sc_hd__buf_6 _7598_ (.A(_2691_),
    .X(_2692_));
 sky130_fd_sc_hd__or2b_2 _7599_ (.A(net127),
    .B_N(_2638_),
    .X(_2693_));
 sky130_fd_sc_hd__nor2_4 _7600_ (.A(net81),
    .B(_2632_),
    .Y(_2694_));
 sky130_fd_sc_hd__nand4_4 _7601_ (.A(net108),
    .B(_2603_),
    .C(_2618_),
    .D(_2596_),
    .Y(_2695_));
 sky130_fd_sc_hd__and4_1 _7602_ (.A(_2616_),
    .B(_2632_),
    .C(_2654_),
    .D(_2695_),
    .X(_2696_));
 sky130_fd_sc_hd__buf_6 _7603_ (.A(_2696_),
    .X(_2697_));
 sky130_fd_sc_hd__o31a_4 _7604_ (.A1(_2659_),
    .A2(_2642_),
    .A3(_2660_),
    .B1(net81),
    .X(_2698_));
 sky130_fd_sc_hd__or4_4 _7605_ (.A(_2693_),
    .B(_2694_),
    .C(_2698_),
    .D(_2697_),
    .X(_2699_));
 sky130_fd_sc_hd__o31ai_4 _7606_ (.A1(_2694_),
    .A2(_2697_),
    .A3(_2698_),
    .B1(_2693_),
    .Y(_2701_));
 sky130_fd_sc_hd__or3b_1 _7607_ (.A(_2598_),
    .B(_2599_),
    .C_N(_2602_),
    .X(_2702_));
 sky130_fd_sc_hd__o21ba_1 _7608_ (.A1(_2672_),
    .A2(_2599_),
    .B1_N(_2598_),
    .X(_2703_));
 sky130_fd_sc_hd__o21a_1 _7609_ (.A1(_2702_),
    .A2(_2666_),
    .B1(_2703_),
    .X(_2704_));
 sky130_fd_sc_hd__nand3_1 _7610_ (.A(_2594_),
    .B(_2618_),
    .C(_2704_),
    .Y(_2705_));
 sky130_fd_sc_hd__nor2_1 _7611_ (.A(net87),
    .B(_2592_),
    .Y(_2706_));
 sky130_fd_sc_hd__o22a_1 _7612_ (.A1(_2706_),
    .A2(_2618_),
    .B1(_2704_),
    .B2(_2596_),
    .X(_2707_));
 sky130_fd_sc_hd__a32oi_4 _7613_ (.A1(_2616_),
    .A2(_2654_),
    .A3(net117),
    .B1(_2705_),
    .B2(_2707_),
    .Y(_2708_));
 sky130_fd_sc_hd__xnor2_2 _7614_ (.A(_2596_),
    .B(_2652_),
    .Y(_2709_));
 sky130_fd_sc_hd__xnor2_2 _7615_ (.A(_2594_),
    .B(_2618_),
    .Y(_2710_));
 sky130_fd_sc_hd__a2111oi_4 _7616_ (.A1(_2709_),
    .A2(_2710_),
    .B1(_2659_),
    .C1(_2660_),
    .D1(_2642_),
    .Y(_2712_));
 sky130_fd_sc_hd__nor2_2 _7617_ (.A(_2708_),
    .B(_2712_),
    .Y(_2713_));
 sky130_fd_sc_hd__and3_1 _7618_ (.A(_2699_),
    .B(_2701_),
    .C(_2713_),
    .X(_2714_));
 sky130_fd_sc_hd__buf_6 _7619_ (.A(_2714_),
    .X(_2715_));
 sky130_fd_sc_hd__buf_6 _7620_ (.A(_2715_),
    .X(_2716_));
 sky130_fd_sc_hd__clkbuf_4 _7621_ (.A(_2633_),
    .X(_2717_));
 sky130_fd_sc_hd__clkbuf_4 _7622_ (.A(_2717_),
    .X(_2718_));
 sky130_fd_sc_hd__or2b_1 _7623_ (.A(net80),
    .B_N(_2718_),
    .X(_2719_));
 sky130_fd_sc_hd__nand3_2 _7624_ (.A(net100),
    .B(_2716_),
    .C(_2719_),
    .Y(_2720_));
 sky130_fd_sc_hd__nor2_1 _7625_ (.A(_2687_),
    .B(_2720_),
    .Y(_2721_));
 sky130_fd_sc_hd__a22o_1 _7626_ (.A1(net80),
    .A2(_2658_),
    .B1(_2680_),
    .B2(_2721_),
    .X(_2723_));
 sky130_fd_sc_hd__clkbuf_4 _7627_ (.A(_2692_),
    .X(_2724_));
 sky130_fd_sc_hd__a32o_2 _7628_ (.A1(_2616_),
    .A2(_2654_),
    .A3(net117),
    .B1(_2705_),
    .B2(_2707_),
    .X(_2725_));
 sky130_fd_sc_hd__a2111o_4 _7629_ (.A1(_2709_),
    .A2(_2710_),
    .B1(_2659_),
    .C1(_2660_),
    .D1(_2642_),
    .X(_2726_));
 sky130_fd_sc_hd__nand2_2 _7630_ (.A(_2725_),
    .B(_2726_),
    .Y(_2727_));
 sky130_fd_sc_hd__buf_2 _7631_ (.A(_2727_),
    .X(_2728_));
 sky130_fd_sc_hd__clkbuf_4 _7632_ (.A(_2633_),
    .X(_2729_));
 sky130_fd_sc_hd__clkbuf_4 _7633_ (.A(_2729_),
    .X(_2730_));
 sky130_fd_sc_hd__a21o_1 _7634_ (.A1(_2533_),
    .A2(_2548_),
    .B1(_2550_),
    .X(_2731_));
 sky130_fd_sc_hd__xnor2_1 _7635_ (.A(_2549_),
    .B(_2551_),
    .Y(_2732_));
 sky130_fd_sc_hd__xnor2_1 _7636_ (.A(_2731_),
    .B(_2732_),
    .Y(_2734_));
 sky130_fd_sc_hd__o31a_1 _7637_ (.A1(_2533_),
    .A2(_2548_),
    .A3(_2552_),
    .B1(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__inv_2 _7638_ (.A(_2735_),
    .Y(_2736_));
 sky130_fd_sc_hd__and2_1 _7639_ (.A(_2730_),
    .B(_2736_),
    .X(_2737_));
 sky130_fd_sc_hd__buf_6 _7640_ (.A(_2699_),
    .X(_2738_));
 sky130_fd_sc_hd__buf_2 _7641_ (.A(_2701_),
    .X(_2739_));
 sky130_fd_sc_hd__and4bb_1 _7642_ (.A_N(_2728_),
    .B_N(_2737_),
    .C(net113),
    .D(_2739_),
    .X(_2740_));
 sky130_fd_sc_hd__nand2_1 _7643_ (.A(_2724_),
    .B(_2740_),
    .Y(_2741_));
 sky130_fd_sc_hd__xnor2_4 _7644_ (.A(net101),
    .B(_2669_),
    .Y(_2742_));
 sky130_fd_sc_hd__nand2_1 _7645_ (.A(net130),
    .B(_2676_),
    .Y(_2743_));
 sky130_fd_sc_hd__or2_1 _7646_ (.A(_2742_),
    .B(_2743_),
    .X(_2745_));
 sky130_fd_sc_hd__buf_2 _7647_ (.A(_2745_),
    .X(_2746_));
 sky130_fd_sc_hd__buf_2 _7648_ (.A(net130),
    .X(_2747_));
 sky130_fd_sc_hd__clkbuf_4 _7649_ (.A(_2747_),
    .X(_2748_));
 sky130_fd_sc_hd__o32a_2 _7650_ (.A1(_2687_),
    .A2(_2741_),
    .A3(_2746_),
    .B1(_2736_),
    .B2(_2748_),
    .X(_2749_));
 sky130_fd_sc_hd__and2_1 _7651_ (.A(_2723_),
    .B(_2749_),
    .X(_2750_));
 sky130_fd_sc_hd__nor2_1 _7652_ (.A(_2723_),
    .B(_2749_),
    .Y(_2751_));
 sky130_fd_sc_hd__nor2_1 _7653_ (.A(_2750_),
    .B(_2751_),
    .Y(_2752_));
 sky130_fd_sc_hd__nand2_1 _7654_ (.A(_2642_),
    .B(_2752_),
    .Y(_2753_));
 sky130_fd_sc_hd__xnor2_4 _7655_ (.A(_2625_),
    .B(_2684_),
    .Y(_2754_));
 sky130_fd_sc_hd__clkbuf_4 _7656_ (.A(_2754_),
    .X(_2756_));
 sky130_fd_sc_hd__buf_2 _7657_ (.A(_2756_),
    .X(_2757_));
 sky130_fd_sc_hd__clkbuf_4 _7658_ (.A(_2692_),
    .X(_2758_));
 sky130_fd_sc_hd__mux2_1 _7659_ (.A0(net79),
    .A1(net78),
    .S(_2730_),
    .X(_2759_));
 sky130_fd_sc_hd__or4_4 _7660_ (.A(_2639_),
    .B(_2694_),
    .C(_2698_),
    .D(_2697_),
    .X(_2760_));
 sky130_fd_sc_hd__o31ai_4 _7661_ (.A1(_2694_),
    .A2(_2697_),
    .A3(_2698_),
    .B1(net107),
    .Y(_2761_));
 sky130_fd_sc_hd__and3_1 _7662_ (.A(_2760_),
    .B(_2761_),
    .C(_2713_),
    .X(_2762_));
 sky130_fd_sc_hd__buf_6 _7663_ (.A(_2762_),
    .X(_2763_));
 sky130_fd_sc_hd__a22o_1 _7664_ (.A1(net132),
    .A2(_2759_),
    .B1(_2763_),
    .B2(_2719_),
    .X(_2764_));
 sky130_fd_sc_hd__and3_1 _7665_ (.A(_2757_),
    .B(_2758_),
    .C(_2764_),
    .X(_2765_));
 sky130_fd_sc_hd__a22o_1 _7666_ (.A1(net78),
    .A2(_2658_),
    .B1(_2680_),
    .B2(_2765_),
    .X(_2767_));
 sky130_fd_sc_hd__nor4_1 _7667_ (.A(_2693_),
    .B(_2694_),
    .C(_2697_),
    .D(_2698_),
    .Y(_2768_));
 sky130_fd_sc_hd__buf_2 _7668_ (.A(_2768_),
    .X(_2769_));
 sky130_fd_sc_hd__o31a_1 _7669_ (.A1(_2694_),
    .A2(_2697_),
    .A3(_2698_),
    .B1(_2693_),
    .X(_2770_));
 sky130_fd_sc_hd__clkbuf_4 _7670_ (.A(_2770_),
    .X(_2771_));
 sky130_fd_sc_hd__and3_1 _7671_ (.A(_0358_),
    .B(_2490_),
    .C(_2512_),
    .X(_2772_));
 sky130_fd_sc_hd__xnor2_1 _7672_ (.A(_2772_),
    .B(_2532_),
    .Y(_2773_));
 sky130_fd_sc_hd__xnor2_1 _7673_ (.A(_2533_),
    .B(_2548_),
    .Y(_2774_));
 sky130_fd_sc_hd__clkbuf_4 _7674_ (.A(_2619_),
    .X(_2775_));
 sky130_fd_sc_hd__mux2_2 _7675_ (.A0(_2773_),
    .A1(_2774_),
    .S(_2775_),
    .X(_2776_));
 sky130_fd_sc_hd__a21oi_1 _7676_ (.A1(_0358_),
    .A2(_2490_),
    .B1(_2512_),
    .Y(_2778_));
 sky130_fd_sc_hd__nor2_1 _7677_ (.A(_2772_),
    .B(_2778_),
    .Y(_2779_));
 sky130_fd_sc_hd__inv_2 _7678_ (.A(_2779_),
    .Y(_2780_));
 sky130_fd_sc_hd__mux2_1 _7679_ (.A0(_2780_),
    .A1(_2773_),
    .S(_2775_),
    .X(_2781_));
 sky130_fd_sc_hd__mux2_1 _7680_ (.A0(_2776_),
    .A1(_2781_),
    .S(_2729_),
    .X(_2782_));
 sky130_fd_sc_hd__or4_1 _7681_ (.A(_2769_),
    .B(_2771_),
    .C(_2727_),
    .D(_2782_),
    .X(_2783_));
 sky130_fd_sc_hd__a211o_1 _7682_ (.A1(net109),
    .A2(_2701_),
    .B1(_2728_),
    .C1(_2737_),
    .X(_2784_));
 sky130_fd_sc_hd__xor2_4 _7683_ (.A(_2629_),
    .B(_2690_),
    .X(_2785_));
 sky130_fd_sc_hd__clkbuf_4 _7684_ (.A(_2785_),
    .X(_2786_));
 sky130_fd_sc_hd__a21oi_1 _7685_ (.A1(_2783_),
    .A2(_2784_),
    .B1(_2786_),
    .Y(_2787_));
 sky130_fd_sc_hd__and4_1 _7686_ (.A(_2747_),
    .B(_2756_),
    .C(_2676_),
    .D(_2787_),
    .X(_2789_));
 sky130_fd_sc_hd__o2bb2a_1 _7687_ (.A1_N(_2670_),
    .A2_N(_2789_),
    .B1(_2781_),
    .B2(_2748_),
    .X(_2790_));
 sky130_fd_sc_hd__nand2_1 _7688_ (.A(_2767_),
    .B(_2790_),
    .Y(_2791_));
 sky130_fd_sc_hd__or2_1 _7689_ (.A(_2767_),
    .B(_2790_),
    .X(_2792_));
 sky130_fd_sc_hd__nand2_2 _7690_ (.A(_2791_),
    .B(_2792_),
    .Y(_2793_));
 sky130_fd_sc_hd__clkbuf_4 _7691_ (.A(_2717_),
    .X(_2794_));
 sky130_fd_sc_hd__a22o_1 _7692_ (.A1(_2699_),
    .A2(_2701_),
    .B1(_2713_),
    .B2(_2794_),
    .X(_2795_));
 sky130_fd_sc_hd__mux2_1 _7693_ (.A0(net80),
    .A1(net79),
    .S(_2633_),
    .X(_2796_));
 sky130_fd_sc_hd__and3_1 _7694_ (.A(_2725_),
    .B(_2726_),
    .C(_2796_),
    .X(_2797_));
 sky130_fd_sc_hd__or3_1 _7695_ (.A(_2769_),
    .B(_2771_),
    .C(_2797_),
    .X(_2798_));
 sky130_fd_sc_hd__and3_1 _7696_ (.A(net100),
    .B(_2795_),
    .C(_2798_),
    .X(_2800_));
 sky130_fd_sc_hd__a32o_1 _7697_ (.A1(_2757_),
    .A2(_2680_),
    .A3(_2800_),
    .B1(_2658_),
    .B2(net79),
    .X(_2801_));
 sky130_fd_sc_hd__clkbuf_4 _7698_ (.A(_2685_),
    .X(_2802_));
 sky130_fd_sc_hd__clkbuf_4 _7699_ (.A(_2692_),
    .X(_2803_));
 sky130_fd_sc_hd__buf_2 _7700_ (.A(_2769_),
    .X(_2804_));
 sky130_fd_sc_hd__buf_2 _7701_ (.A(_2771_),
    .X(_2805_));
 sky130_fd_sc_hd__mux2_1 _7702_ (.A0(_2736_),
    .A1(_2776_),
    .S(_2717_),
    .X(_2806_));
 sky130_fd_sc_hd__nor3_1 _7703_ (.A(_2708_),
    .B(_2712_),
    .C(_2806_),
    .Y(_2807_));
 sky130_fd_sc_hd__or3_1 _7704_ (.A(_2804_),
    .B(_2805_),
    .C(_2807_),
    .X(_2808_));
 sky130_fd_sc_hd__nand3_1 _7705_ (.A(_2803_),
    .B(_2795_),
    .C(_2808_),
    .Y(_2809_));
 sky130_fd_sc_hd__or3_1 _7706_ (.A(_2802_),
    .B(_2743_),
    .C(_2809_),
    .X(_2811_));
 sky130_fd_sc_hd__clkbuf_4 _7707_ (.A(_2742_),
    .X(_2812_));
 sky130_fd_sc_hd__o22a_1 _7708_ (.A1(_2748_),
    .A2(_2776_),
    .B1(_2811_),
    .B2(_2812_),
    .X(_2813_));
 sky130_fd_sc_hd__nor2_1 _7709_ (.A(_2801_),
    .B(_2813_),
    .Y(_2814_));
 sky130_fd_sc_hd__nand2_1 _7710_ (.A(_2801_),
    .B(_2813_),
    .Y(_2815_));
 sky130_fd_sc_hd__nand2b_2 _7711_ (.A_N(_2814_),
    .B(_2815_),
    .Y(_2816_));
 sky130_fd_sc_hd__or2_1 _7712_ (.A(_2793_),
    .B(_2816_),
    .X(_2817_));
 sky130_fd_sc_hd__or2_2 _7713_ (.A(_2753_),
    .B(_2817_),
    .X(_2818_));
 sky130_fd_sc_hd__and2_2 _7714_ (.A(_2661_),
    .B(_2676_),
    .X(_2819_));
 sky130_fd_sc_hd__nand2_1 _7715_ (.A(_2670_),
    .B(_2819_),
    .Y(_2820_));
 sky130_fd_sc_hd__a21o_1 _7716_ (.A1(_2794_),
    .A2(_2716_),
    .B1(_2724_),
    .X(_2822_));
 sky130_fd_sc_hd__nand2_4 _7717_ (.A(_2699_),
    .B(_2701_),
    .Y(_2823_));
 sky130_fd_sc_hd__clkbuf_4 _7718_ (.A(_2823_),
    .X(_2824_));
 sky130_fd_sc_hd__mux2_1 _7719_ (.A0(net78),
    .A1(net76),
    .S(_2729_),
    .X(_2825_));
 sky130_fd_sc_hd__a221o_1 _7720_ (.A1(_2824_),
    .A2(_2797_),
    .B1(_2716_),
    .B2(_2825_),
    .C1(_2786_),
    .X(_2826_));
 sky130_fd_sc_hd__nand2_1 _7721_ (.A(_2822_),
    .B(_2826_),
    .Y(_2827_));
 sky130_fd_sc_hd__inv_2 _7722_ (.A(net76),
    .Y(_2828_));
 sky130_fd_sc_hd__o32a_1 _7723_ (.A1(_2687_),
    .A2(_2820_),
    .A3(_2827_),
    .B1(_2661_),
    .B2(_2828_),
    .X(_2829_));
 sky130_fd_sc_hd__nor2_2 _7724_ (.A(_2655_),
    .B(_2642_),
    .Y(_2830_));
 sky130_fd_sc_hd__clkbuf_4 _7725_ (.A(_2830_),
    .X(_2831_));
 sky130_fd_sc_hd__xor2_1 _7726_ (.A(_0358_),
    .B(_2490_),
    .X(_2833_));
 sky130_fd_sc_hd__mux2_1 _7727_ (.A0(_2833_),
    .A1(_2779_),
    .S(_2619_),
    .X(_2834_));
 sky130_fd_sc_hd__clkbuf_4 _7728_ (.A(_2756_),
    .X(_2835_));
 sky130_fd_sc_hd__inv_2 _7729_ (.A(_2834_),
    .Y(_2836_));
 sky130_fd_sc_hd__mux2_1 _7730_ (.A0(_2781_),
    .A1(_2836_),
    .S(_2729_),
    .X(_2837_));
 sky130_fd_sc_hd__or4_1 _7731_ (.A(_2769_),
    .B(_2771_),
    .C(_2727_),
    .D(_2837_),
    .X(_2838_));
 sky130_fd_sc_hd__o21ai_1 _7732_ (.A1(_2769_),
    .A2(_2771_),
    .B1(_2807_),
    .Y(_2839_));
 sky130_fd_sc_hd__nand3_1 _7733_ (.A(_2758_),
    .B(_2838_),
    .C(_2839_),
    .Y(_2840_));
 sky130_fd_sc_hd__and3_1 _7734_ (.A(_2835_),
    .B(_2822_),
    .C(_2840_),
    .X(_2841_));
 sky130_fd_sc_hd__and3_1 _7735_ (.A(net130),
    .B(_2670_),
    .C(_2676_),
    .X(_2842_));
 sky130_fd_sc_hd__clkbuf_4 _7736_ (.A(_2842_),
    .X(_2844_));
 sky130_fd_sc_hd__a22o_1 _7737_ (.A1(_2831_),
    .A2(_2834_),
    .B1(_2841_),
    .B2(_2844_),
    .X(_2845_));
 sky130_fd_sc_hd__or2_1 _7738_ (.A(_2829_),
    .B(_2845_),
    .X(_2846_));
 sky130_fd_sc_hd__nand2_1 _7739_ (.A(_2829_),
    .B(_2845_),
    .Y(_2847_));
 sky130_fd_sc_hd__nand2_2 _7740_ (.A(_2846_),
    .B(_2847_),
    .Y(_2848_));
 sky130_fd_sc_hd__a21o_1 _7741_ (.A1(_2716_),
    .A2(_2719_),
    .B1(_2724_),
    .X(_2849_));
 sky130_fd_sc_hd__buf_2 _7742_ (.A(_2725_),
    .X(_2850_));
 sky130_fd_sc_hd__buf_2 _7743_ (.A(_2726_),
    .X(_2851_));
 sky130_fd_sc_hd__mux2_1 _7744_ (.A0(net76),
    .A1(net75),
    .S(_2729_),
    .X(_2852_));
 sky130_fd_sc_hd__and3_1 _7745_ (.A(_2850_),
    .B(_2851_),
    .C(_2852_),
    .X(_2853_));
 sky130_fd_sc_hd__nor2_2 _7746_ (.A(_2768_),
    .B(_2770_),
    .Y(_2855_));
 sky130_fd_sc_hd__clkbuf_4 _7747_ (.A(_2855_),
    .X(_2856_));
 sky130_fd_sc_hd__a221o_1 _7748_ (.A1(_2759_),
    .A2(_2763_),
    .B1(_2853_),
    .B2(_2856_),
    .C1(_2786_),
    .X(_2857_));
 sky130_fd_sc_hd__and3_1 _7749_ (.A(_2757_),
    .B(_2849_),
    .C(_2857_),
    .X(_2858_));
 sky130_fd_sc_hd__a22o_1 _7750_ (.A1(net75),
    .A2(_2658_),
    .B1(_2680_),
    .B2(_2858_),
    .X(_2859_));
 sky130_fd_sc_hd__or2_1 _7751_ (.A(_2724_),
    .B(_2740_),
    .X(_2860_));
 sky130_fd_sc_hd__a211oi_1 _7752_ (.A1(_2699_),
    .A2(_2701_),
    .B1(_2727_),
    .C1(_2782_),
    .Y(_2861_));
 sky130_fd_sc_hd__nor3_1 _7753_ (.A(_2328_),
    .B(_2349_),
    .C(_2486_),
    .Y(_2862_));
 sky130_fd_sc_hd__and2b_1 _7754_ (.A_N(_2862_),
    .B(_2487_),
    .X(_2863_));
 sky130_fd_sc_hd__nor2_1 _7755_ (.A(_2489_),
    .B(_2863_),
    .Y(_2864_));
 sky130_fd_sc_hd__or2_1 _7756_ (.A(_2490_),
    .B(_2864_),
    .X(_2866_));
 sky130_fd_sc_hd__inv_2 _7757_ (.A(_2833_),
    .Y(_2867_));
 sky130_fd_sc_hd__mux2_1 _7758_ (.A0(_2866_),
    .A1(_2867_),
    .S(_2775_),
    .X(_2868_));
 sky130_fd_sc_hd__mux2_1 _7759_ (.A0(_2836_),
    .A1(_2868_),
    .S(_2717_),
    .X(_2869_));
 sky130_fd_sc_hd__a211oi_1 _7760_ (.A1(net125),
    .A2(_2761_),
    .B1(_2727_),
    .C1(_2869_),
    .Y(_2870_));
 sky130_fd_sc_hd__or3_1 _7761_ (.A(_2786_),
    .B(_2861_),
    .C(_2870_),
    .X(_2871_));
 sky130_fd_sc_hd__nand2_1 _7762_ (.A(_2860_),
    .B(_2871_),
    .Y(_2872_));
 sky130_fd_sc_hd__o32a_1 _7763_ (.A1(_2687_),
    .A2(_2746_),
    .A3(_2872_),
    .B1(_2868_),
    .B2(_2747_),
    .X(_2873_));
 sky130_fd_sc_hd__nand2_1 _7764_ (.A(_2859_),
    .B(_2873_),
    .Y(_2874_));
 sky130_fd_sc_hd__or2_1 _7765_ (.A(_2859_),
    .B(_2873_),
    .X(_2875_));
 sky130_fd_sc_hd__nand2_2 _7766_ (.A(_2874_),
    .B(_2875_),
    .Y(_2877_));
 sky130_fd_sc_hd__nor2_1 _7767_ (.A(_2848_),
    .B(_2877_),
    .Y(_2878_));
 sky130_fd_sc_hd__a21o_1 _7768_ (.A1(_2795_),
    .A2(_2808_),
    .B1(_2803_),
    .X(_2879_));
 sky130_fd_sc_hd__clkbuf_4 _7769_ (.A(_2785_),
    .X(_2880_));
 sky130_fd_sc_hd__and4b_1 _7770_ (.A_N(_2837_),
    .B(_2761_),
    .C(net125),
    .D(_2713_),
    .X(_2881_));
 sky130_fd_sc_hd__and2b_1 _7771_ (.A_N(_2487_),
    .B(_2862_),
    .X(_2882_));
 sky130_fd_sc_hd__nor2_1 _7772_ (.A(_2863_),
    .B(_2882_),
    .Y(_2883_));
 sky130_fd_sc_hd__inv_2 _7773_ (.A(_2866_),
    .Y(_2884_));
 sky130_fd_sc_hd__mux2_1 _7774_ (.A0(_2883_),
    .A1(_2884_),
    .S(_2619_),
    .X(_2885_));
 sky130_fd_sc_hd__inv_2 _7775_ (.A(_2885_),
    .Y(_2886_));
 sky130_fd_sc_hd__mux2_1 _7776_ (.A0(_2868_),
    .A1(_2886_),
    .S(_2729_),
    .X(_2888_));
 sky130_fd_sc_hd__or3_1 _7777_ (.A(_2708_),
    .B(_2712_),
    .C(_2888_),
    .X(_2889_));
 sky130_fd_sc_hd__a21oi_1 _7778_ (.A1(net122),
    .A2(_2761_),
    .B1(_2889_),
    .Y(_2890_));
 sky130_fd_sc_hd__or3_4 _7779_ (.A(_2880_),
    .B(_2881_),
    .C(_2890_),
    .X(_2891_));
 sky130_fd_sc_hd__nor2_1 _7780_ (.A(_2747_),
    .B(_2886_),
    .Y(_2892_));
 sky130_fd_sc_hd__a41o_1 _7781_ (.A1(_2757_),
    .A2(_2844_),
    .A3(_2879_),
    .A4(_2891_),
    .B1(_2892_),
    .X(_2893_));
 sky130_fd_sc_hd__a21o_1 _7782_ (.A1(_2795_),
    .A2(_2798_),
    .B1(_2803_),
    .X(_2894_));
 sky130_fd_sc_hd__buf_6 _7783_ (.A(_2763_),
    .X(_2895_));
 sky130_fd_sc_hd__mux2_1 _7784_ (.A0(net75),
    .A1(net74),
    .S(_2633_),
    .X(_2896_));
 sky130_fd_sc_hd__and3_1 _7785_ (.A(_2850_),
    .B(_2851_),
    .C(_2896_),
    .X(_2897_));
 sky130_fd_sc_hd__a221o_1 _7786_ (.A1(_2895_),
    .A2(_2825_),
    .B1(_2897_),
    .B2(_2856_),
    .C1(_2880_),
    .X(_2899_));
 sky130_fd_sc_hd__and3_1 _7787_ (.A(_2757_),
    .B(_2894_),
    .C(_2899_),
    .X(_2900_));
 sky130_fd_sc_hd__a22o_1 _7788_ (.A1(net74),
    .A2(_2658_),
    .B1(_2680_),
    .B2(_2900_),
    .X(_2901_));
 sky130_fd_sc_hd__and2b_1 _7789_ (.A_N(_2893_),
    .B(_2901_),
    .X(_2902_));
 sky130_fd_sc_hd__or2b_1 _7790_ (.A(_2901_),
    .B_N(_2893_),
    .X(_2903_));
 sky130_fd_sc_hd__nand2b_2 _7791_ (.A_N(_2902_),
    .B(_2903_),
    .Y(_2904_));
 sky130_fd_sc_hd__or2_1 _7792_ (.A(_2355_),
    .B(_2479_),
    .X(_2905_));
 sky130_fd_sc_hd__and2b_1 _7793_ (.A_N(_2905_),
    .B(_2481_),
    .X(_2906_));
 sky130_fd_sc_hd__nor2_1 _7794_ (.A(_2346_),
    .B(_2906_),
    .Y(_2907_));
 sky130_fd_sc_hd__o21ba_1 _7795_ (.A1(_2342_),
    .A2(_2907_),
    .B1_N(_2347_),
    .X(_2908_));
 sky130_fd_sc_hd__o21ai_1 _7796_ (.A1(_2336_),
    .A2(_2908_),
    .B1(_2484_),
    .Y(_2910_));
 sky130_fd_sc_hd__xnor2_1 _7797_ (.A(_2331_),
    .B(_2910_),
    .Y(_2911_));
 sky130_fd_sc_hd__mux2_1 _7798_ (.A0(_2911_),
    .A1(_2883_),
    .S(_2619_),
    .X(_2912_));
 sky130_fd_sc_hd__clkbuf_4 _7799_ (.A(_2880_),
    .X(_2913_));
 sky130_fd_sc_hd__nand3_1 _7800_ (.A(_2913_),
    .B(_2783_),
    .C(_2784_),
    .Y(_2914_));
 sky130_fd_sc_hd__nor2_1 _7801_ (.A(_2727_),
    .B(_2869_),
    .Y(_2915_));
 sky130_fd_sc_hd__mux2_1 _7802_ (.A0(_2885_),
    .A1(_2912_),
    .S(_2633_),
    .X(_2916_));
 sky130_fd_sc_hd__buf_6 _7803_ (.A(_2715_),
    .X(_2917_));
 sky130_fd_sc_hd__clkbuf_4 _7804_ (.A(_2785_),
    .X(_2918_));
 sky130_fd_sc_hd__a221o_1 _7805_ (.A1(_2824_),
    .A2(_2915_),
    .B1(_2916_),
    .B2(_2917_),
    .C1(_2918_),
    .X(_2919_));
 sky130_fd_sc_hd__and3_1 _7806_ (.A(_2757_),
    .B(_2914_),
    .C(_2919_),
    .X(_2921_));
 sky130_fd_sc_hd__a22o_1 _7807_ (.A1(_2831_),
    .A2(_2912_),
    .B1(_2921_),
    .B2(_2844_),
    .X(_2922_));
 sky130_fd_sc_hd__clkbuf_4 _7808_ (.A(_2754_),
    .X(_2923_));
 sky130_fd_sc_hd__a221o_1 _7809_ (.A1(_2716_),
    .A2(_2759_),
    .B1(_2895_),
    .B2(_2719_),
    .C1(_2724_),
    .X(_2924_));
 sky130_fd_sc_hd__mux2_1 _7810_ (.A0(net74),
    .A1(net73),
    .S(_2730_),
    .X(_2925_));
 sky130_fd_sc_hd__a221o_1 _7811_ (.A1(_2824_),
    .A2(_2853_),
    .B1(_2925_),
    .B2(_2716_),
    .C1(_2880_),
    .X(_2926_));
 sky130_fd_sc_hd__and4_1 _7812_ (.A(_2926_),
    .B(_2819_),
    .C(_2924_),
    .D(_2923_),
    .X(_2927_));
 sky130_fd_sc_hd__a22o_1 _7813_ (.A1(net73),
    .A2(_2658_),
    .B1(_2670_),
    .B2(_2927_),
    .X(_2928_));
 sky130_fd_sc_hd__or2b_1 _7814_ (.A(_2922_),
    .B_N(_2928_),
    .X(_2929_));
 sky130_fd_sc_hd__or2b_1 _7815_ (.A(_2928_),
    .B_N(_2922_),
    .X(_2930_));
 sky130_fd_sc_hd__nand2_2 _7816_ (.A(_2929_),
    .B(_2930_),
    .Y(_2932_));
 sky130_fd_sc_hd__nor2_1 _7817_ (.A(_2904_),
    .B(_2932_),
    .Y(_2933_));
 sky130_fd_sc_hd__and2_1 _7818_ (.A(_2878_),
    .B(_2933_),
    .X(_2934_));
 sky130_fd_sc_hd__mux2_1 _7819_ (.A0(net96),
    .A1(net95),
    .S(_2730_),
    .X(_2935_));
 sky130_fd_sc_hd__mux2_1 _7820_ (.A0(net67),
    .A1(net97),
    .S(_2717_),
    .X(_2936_));
 sky130_fd_sc_hd__and3_1 _7821_ (.A(_2850_),
    .B(_2851_),
    .C(_2936_),
    .X(_2937_));
 sky130_fd_sc_hd__a22o_1 _7822_ (.A1(_2715_),
    .A2(_2935_),
    .B1(_2937_),
    .B2(_2823_),
    .X(_2938_));
 sky130_fd_sc_hd__mux2_1 _7823_ (.A0(net69),
    .A1(net68),
    .S(_2717_),
    .X(_2939_));
 sky130_fd_sc_hd__mux2_1 _7824_ (.A0(net71),
    .A1(net70),
    .S(_2729_),
    .X(_2940_));
 sky130_fd_sc_hd__and3_1 _7825_ (.A(_2850_),
    .B(_2851_),
    .C(_2940_),
    .X(_2941_));
 sky130_fd_sc_hd__a22o_1 _7826_ (.A1(_2715_),
    .A2(_2939_),
    .B1(_2941_),
    .B2(_2823_),
    .X(_2943_));
 sky130_fd_sc_hd__mux2_1 _7827_ (.A0(_2938_),
    .A1(_2943_),
    .S(_2880_),
    .X(_2944_));
 sky130_fd_sc_hd__a221o_1 _7828_ (.A1(_2823_),
    .A2(_2797_),
    .B1(_2825_),
    .B2(net132),
    .C1(net100),
    .X(_2945_));
 sky130_fd_sc_hd__mux2_1 _7829_ (.A0(net73),
    .A1(net72),
    .S(_2729_),
    .X(_2946_));
 sky130_fd_sc_hd__a221o_1 _7830_ (.A1(_2823_),
    .A2(_2897_),
    .B1(_2946_),
    .B2(_2715_),
    .C1(_2785_),
    .X(_2947_));
 sky130_fd_sc_hd__and3_1 _7831_ (.A(_2686_),
    .B(_2945_),
    .C(_2947_),
    .X(_2948_));
 sky130_fd_sc_hd__a211o_1 _7832_ (.A1(_2835_),
    .A2(_2944_),
    .B1(_2948_),
    .C1(_2812_),
    .X(_2949_));
 sky130_fd_sc_hd__a41o_1 _7833_ (.A1(_2794_),
    .A2(_2754_),
    .A3(_2803_),
    .A4(_2917_),
    .B1(_2670_),
    .X(_2950_));
 sky130_fd_sc_hd__nand2_1 _7834_ (.A(_2676_),
    .B(_2950_),
    .Y(_2951_));
 sky130_fd_sc_hd__nor2_1 _7835_ (.A(_2657_),
    .B(_2951_),
    .Y(_2952_));
 sky130_fd_sc_hd__a22o_4 _7836_ (.A1(net95),
    .A2(_2657_),
    .B1(_2949_),
    .B2(_2952_),
    .X(_2954_));
 sky130_fd_sc_hd__nor2_1 _7837_ (.A(_2468_),
    .B(_2361_),
    .Y(_2955_));
 sky130_fd_sc_hd__xor2_1 _7838_ (.A(_2955_),
    .B(_2467_),
    .X(_2956_));
 sky130_fd_sc_hd__xnor2_1 _7839_ (.A(_2470_),
    .B(_2475_),
    .Y(_2957_));
 sky130_fd_sc_hd__clkbuf_4 _7840_ (.A(_2619_),
    .X(_2958_));
 sky130_fd_sc_hd__mux2_1 _7841_ (.A0(_2956_),
    .A1(_2957_),
    .S(_2958_),
    .X(_2959_));
 sky130_fd_sc_hd__xnor2_1 _7842_ (.A(_2460_),
    .B(_2465_),
    .Y(_2960_));
 sky130_fd_sc_hd__mux2_1 _7843_ (.A0(_2960_),
    .A1(_2956_),
    .S(_2958_),
    .X(_2961_));
 sky130_fd_sc_hd__or2b_1 _7844_ (.A(_2961_),
    .B_N(_2718_),
    .X(_2962_));
 sky130_fd_sc_hd__o21ai_1 _7845_ (.A1(_2794_),
    .A2(_2959_),
    .B1(_2962_),
    .Y(_2963_));
 sky130_fd_sc_hd__xor2_1 _7846_ (.A(_2368_),
    .B(_2459_),
    .X(_2965_));
 sky130_fd_sc_hd__nand2_1 _7847_ (.A(_2775_),
    .B(_2960_),
    .Y(_2966_));
 sky130_fd_sc_hd__o21ai_2 _7848_ (.A1(_2775_),
    .A2(_2965_),
    .B1(_2966_),
    .Y(_2967_));
 sky130_fd_sc_hd__inv_2 _7849_ (.A(_2967_),
    .Y(_2968_));
 sky130_fd_sc_hd__xor2_1 _7850_ (.A(_2374_),
    .B(_2456_),
    .X(_2969_));
 sky130_fd_sc_hd__mux2_1 _7851_ (.A0(_2969_),
    .A1(_2965_),
    .S(_2775_),
    .X(_2970_));
 sky130_fd_sc_hd__mux2_1 _7852_ (.A0(_2968_),
    .A1(_2970_),
    .S(_2717_),
    .X(_2971_));
 sky130_fd_sc_hd__or3b_1 _7853_ (.A(_2708_),
    .B(_2712_),
    .C_N(_2971_),
    .X(_2972_));
 sky130_fd_sc_hd__o2bb2a_1 _7854_ (.A1_N(_2763_),
    .A2_N(_2963_),
    .B1(_2972_),
    .B2(_2823_),
    .X(_2973_));
 sky130_fd_sc_hd__xnor2_1 _7855_ (.A(_2482_),
    .B(_2907_),
    .Y(_2974_));
 sky130_fd_sc_hd__xor2_1 _7856_ (.A(_2336_),
    .B(_2908_),
    .X(_2976_));
 sky130_fd_sc_hd__mux2_2 _7857_ (.A0(_2974_),
    .A1(_2976_),
    .S(_2619_),
    .X(_2977_));
 sky130_fd_sc_hd__and2b_1 _7858_ (.A_N(_2481_),
    .B(_2905_),
    .X(_2978_));
 sky130_fd_sc_hd__or2_1 _7859_ (.A(_2906_),
    .B(_2978_),
    .X(_2979_));
 sky130_fd_sc_hd__nor2_1 _7860_ (.A(_2775_),
    .B(_2979_),
    .Y(_2980_));
 sky130_fd_sc_hd__a21oi_2 _7861_ (.A1(_2775_),
    .A2(_2974_),
    .B1(_2980_),
    .Y(_2981_));
 sky130_fd_sc_hd__inv_2 _7862_ (.A(_2981_),
    .Y(_2982_));
 sky130_fd_sc_hd__mux2_1 _7863_ (.A0(_2977_),
    .A1(_2982_),
    .S(_2717_),
    .X(_2983_));
 sky130_fd_sc_hd__o21ai_1 _7864_ (.A1(_2470_),
    .A2(_2475_),
    .B1(_2478_),
    .Y(_2984_));
 sky130_fd_sc_hd__or2_1 _7865_ (.A(_2476_),
    .B(_2355_),
    .X(_2985_));
 sky130_fd_sc_hd__xnor2_1 _7866_ (.A(_2984_),
    .B(_2985_),
    .Y(_2987_));
 sky130_fd_sc_hd__nor2_1 _7867_ (.A(_2775_),
    .B(_2987_),
    .Y(_2988_));
 sky130_fd_sc_hd__a21oi_1 _7868_ (.A1(_2958_),
    .A2(_2979_),
    .B1(_2988_),
    .Y(_2989_));
 sky130_fd_sc_hd__inv_2 _7869_ (.A(_2989_),
    .Y(_2990_));
 sky130_fd_sc_hd__inv_2 _7870_ (.A(_2987_),
    .Y(_2991_));
 sky130_fd_sc_hd__mux2_1 _7871_ (.A0(_2957_),
    .A1(_2991_),
    .S(_2958_),
    .X(_2992_));
 sky130_fd_sc_hd__mux2_1 _7872_ (.A0(_2990_),
    .A1(_2992_),
    .S(_2717_),
    .X(_2993_));
 sky130_fd_sc_hd__or2_1 _7873_ (.A(_2728_),
    .B(_2993_),
    .X(_2994_));
 sky130_fd_sc_hd__o2bb2a_1 _7874_ (.A1_N(_2763_),
    .A2_N(_2983_),
    .B1(_2994_),
    .B2(_2823_),
    .X(_2995_));
 sky130_fd_sc_hd__mux2_1 _7875_ (.A0(_2973_),
    .A1(_2995_),
    .S(_2918_),
    .X(_2996_));
 sky130_fd_sc_hd__and3_1 _7876_ (.A(_2785_),
    .B(_2838_),
    .C(_2839_),
    .X(_2998_));
 sky130_fd_sc_hd__mux2_1 _7877_ (.A0(_2976_),
    .A1(_2911_),
    .S(_2619_),
    .X(_2999_));
 sky130_fd_sc_hd__mux2_1 _7878_ (.A0(_2912_),
    .A1(_2999_),
    .S(_2633_),
    .X(_3000_));
 sky130_fd_sc_hd__and3_1 _7879_ (.A(_2725_),
    .B(_2726_),
    .C(_3000_),
    .X(_3001_));
 sky130_fd_sc_hd__or3_1 _7880_ (.A(_2769_),
    .B(_2771_),
    .C(_3001_),
    .X(_3002_));
 sky130_fd_sc_hd__o21ai_1 _7881_ (.A1(_2804_),
    .A2(_2805_),
    .B1(_2889_),
    .Y(_3003_));
 sky130_fd_sc_hd__a21oi_1 _7882_ (.A1(_3002_),
    .A2(_3003_),
    .B1(_2880_),
    .Y(_3004_));
 sky130_fd_sc_hd__o31a_1 _7883_ (.A1(_2756_),
    .A2(_2998_),
    .A3(_3004_),
    .B1(_2670_),
    .X(_3005_));
 sky130_fd_sc_hd__o21a_1 _7884_ (.A1(_2687_),
    .A2(_2996_),
    .B1(_3005_),
    .X(_3006_));
 sky130_fd_sc_hd__nand2_1 _7885_ (.A(_2831_),
    .B(_2970_),
    .Y(_3007_));
 sky130_fd_sc_hd__o31a_2 _7886_ (.A1(_2831_),
    .A2(_2951_),
    .A3(_3006_),
    .B1(_3007_),
    .X(_3009_));
 sky130_fd_sc_hd__xor2_4 _7887_ (.A(_2954_),
    .B(_3009_),
    .X(_3010_));
 sky130_fd_sc_hd__mux2_2 _7888_ (.A0(net70),
    .A1(net69),
    .S(_2730_),
    .X(_3011_));
 sky130_fd_sc_hd__mux2_1 _7889_ (.A0(net68),
    .A1(net67),
    .S(_2718_),
    .X(_3012_));
 sky130_fd_sc_hd__a22o_1 _7890_ (.A1(_2895_),
    .A2(_3011_),
    .B1(_3012_),
    .B2(_2917_),
    .X(_3013_));
 sky130_fd_sc_hd__buf_2 _7891_ (.A(_2713_),
    .X(_3014_));
 sky130_fd_sc_hd__mux2_1 _7892_ (.A0(net97),
    .A1(net96),
    .S(_2730_),
    .X(_3015_));
 sky130_fd_sc_hd__o211a_1 _7893_ (.A1(_2804_),
    .A2(_2805_),
    .B1(_3014_),
    .C1(_3015_),
    .X(_3016_));
 sky130_fd_sc_hd__mux2_1 _7894_ (.A0(net95),
    .A1(net94),
    .S(_2718_),
    .X(_3017_));
 sky130_fd_sc_hd__and4_1 _7895_ (.A(net113),
    .B(_2739_),
    .C(_3014_),
    .D(_3017_),
    .X(_3018_));
 sky130_fd_sc_hd__o21a_1 _7896_ (.A1(_3016_),
    .A2(_3018_),
    .B1(_2803_),
    .X(_3020_));
 sky130_fd_sc_hd__a211o_1 _7897_ (.A1(_2913_),
    .A2(_3013_),
    .B1(_3020_),
    .C1(_2802_),
    .X(_3021_));
 sky130_fd_sc_hd__a221o_1 _7898_ (.A1(_2759_),
    .A2(_2763_),
    .B1(_2853_),
    .B2(_2856_),
    .C1(net100),
    .X(_3022_));
 sky130_fd_sc_hd__mux2_1 _7899_ (.A0(net72),
    .A1(net71),
    .S(_2730_),
    .X(_3023_));
 sky130_fd_sc_hd__a221o_1 _7900_ (.A1(_2763_),
    .A2(_2925_),
    .B1(_3023_),
    .B2(net106),
    .C1(_2785_),
    .X(_3024_));
 sky130_fd_sc_hd__a21o_1 _7901_ (.A1(_3022_),
    .A2(_3024_),
    .B1(_2923_),
    .X(_3025_));
 sky130_fd_sc_hd__a21o_1 _7902_ (.A1(_3021_),
    .A2(_3025_),
    .B1(_2812_),
    .X(_3026_));
 sky130_fd_sc_hd__nand2_1 _7903_ (.A(_2835_),
    .B(_2819_),
    .Y(_3027_));
 sky130_fd_sc_hd__o21ai_2 _7904_ (.A1(_3027_),
    .A2(_2720_),
    .B1(_2820_),
    .Y(_3028_));
 sky130_fd_sc_hd__a22oi_4 _7905_ (.A1(net94),
    .A2(_2657_),
    .B1(_3026_),
    .B2(_3028_),
    .Y(_3029_));
 sky130_fd_sc_hd__or2b_1 _7906_ (.A(_2455_),
    .B_N(_2380_),
    .X(_3031_));
 sky130_fd_sc_hd__xnor2_1 _7907_ (.A(_3031_),
    .B(_2454_),
    .Y(_3032_));
 sky130_fd_sc_hd__mux2_1 _7908_ (.A0(_3032_),
    .A1(_2969_),
    .S(_2775_),
    .X(_3033_));
 sky130_fd_sc_hd__clkbuf_4 _7909_ (.A(_2686_),
    .X(_3034_));
 sky130_fd_sc_hd__o31a_1 _7910_ (.A1(_3034_),
    .A2(_2743_),
    .A3(_2741_),
    .B1(_2746_),
    .X(_3035_));
 sky130_fd_sc_hd__mux2_1 _7911_ (.A0(_2992_),
    .A1(_2959_),
    .S(_2718_),
    .X(_3036_));
 sky130_fd_sc_hd__inv_2 _7912_ (.A(_3036_),
    .Y(_3037_));
 sky130_fd_sc_hd__nand2_1 _7913_ (.A(_2730_),
    .B(_2990_),
    .Y(_3038_));
 sky130_fd_sc_hd__o211a_1 _7914_ (.A1(_2730_),
    .A2(_2982_),
    .B1(_3038_),
    .C1(_2713_),
    .X(_3039_));
 sky130_fd_sc_hd__a22o_1 _7915_ (.A1(_2917_),
    .A2(_3037_),
    .B1(_3039_),
    .B2(_2824_),
    .X(_3040_));
 sky130_fd_sc_hd__mux2_1 _7916_ (.A0(_2961_),
    .A1(_2967_),
    .S(_2718_),
    .X(_3042_));
 sky130_fd_sc_hd__nor2_1 _7917_ (.A(_2728_),
    .B(_3042_),
    .Y(_3043_));
 sky130_fd_sc_hd__mux2_1 _7918_ (.A0(_2970_),
    .A1(_3033_),
    .S(_2729_),
    .X(_3044_));
 sky130_fd_sc_hd__and3_1 _7919_ (.A(_2850_),
    .B(_2851_),
    .C(_3044_),
    .X(_3045_));
 sky130_fd_sc_hd__or3_1 _7920_ (.A(_2804_),
    .B(_2771_),
    .C(_3045_),
    .X(_3046_));
 sky130_fd_sc_hd__o211a_1 _7921_ (.A1(_2856_),
    .A2(_3043_),
    .B1(_3046_),
    .C1(_2803_),
    .X(_3047_));
 sky130_fd_sc_hd__a21o_1 _7922_ (.A1(_2913_),
    .A2(_3040_),
    .B1(_3047_),
    .X(_3048_));
 sky130_fd_sc_hd__or3_1 _7923_ (.A(_2691_),
    .B(_2861_),
    .C(_2870_),
    .X(_3049_));
 sky130_fd_sc_hd__mux2_1 _7924_ (.A0(_2999_),
    .A1(_2977_),
    .S(_2633_),
    .X(_3050_));
 sky130_fd_sc_hd__and3_1 _7925_ (.A(_2725_),
    .B(_2726_),
    .C(_3050_),
    .X(_3051_));
 sky130_fd_sc_hd__or3_1 _7926_ (.A(_2769_),
    .B(_2771_),
    .C(_3051_),
    .X(_3053_));
 sky130_fd_sc_hd__and3_1 _7927_ (.A(_2725_),
    .B(_2726_),
    .C(_2916_),
    .X(_3054_));
 sky130_fd_sc_hd__a21o_1 _7928_ (.A1(_2699_),
    .A2(_2701_),
    .B1(_3054_),
    .X(_3055_));
 sky130_fd_sc_hd__a21o_1 _7929_ (.A1(_3053_),
    .A2(_3055_),
    .B1(_2785_),
    .X(_3056_));
 sky130_fd_sc_hd__and3_1 _7930_ (.A(_2802_),
    .B(_3049_),
    .C(_3056_),
    .X(_3057_));
 sky130_fd_sc_hd__a211oi_1 _7931_ (.A1(_2757_),
    .A2(_3048_),
    .B1(_3057_),
    .C1(_2812_),
    .Y(_3058_));
 sky130_fd_sc_hd__o2bb2a_2 _7932_ (.A1_N(_2831_),
    .A2_N(_3033_),
    .B1(_3035_),
    .B2(_3058_),
    .X(_3059_));
 sky130_fd_sc_hd__xnor2_4 _7933_ (.A(_3029_),
    .B(_3059_),
    .Y(_3060_));
 sky130_fd_sc_hd__nand2_1 _7934_ (.A(net92),
    .B(_2657_),
    .Y(_3061_));
 sky130_fd_sc_hd__o211a_1 _7935_ (.A1(_2804_),
    .A2(_2805_),
    .B1(_3014_),
    .C1(_3017_),
    .X(_3062_));
 sky130_fd_sc_hd__mux2_1 _7936_ (.A0(net93),
    .A1(net92),
    .S(_2718_),
    .X(_3064_));
 sky130_fd_sc_hd__and4_1 _7937_ (.A(_2738_),
    .B(_2739_),
    .C(_3014_),
    .D(_3064_),
    .X(_3065_));
 sky130_fd_sc_hd__o21ai_1 _7938_ (.A1(_3062_),
    .A2(_3065_),
    .B1(_2758_),
    .Y(_3066_));
 sky130_fd_sc_hd__o211a_1 _7939_ (.A1(_2804_),
    .A2(_2805_),
    .B1(_3014_),
    .C1(_3012_),
    .X(_3067_));
 sky130_fd_sc_hd__and4_1 _7940_ (.A(_2738_),
    .B(_2739_),
    .C(_2713_),
    .D(_3015_),
    .X(_3068_));
 sky130_fd_sc_hd__o21ai_1 _7941_ (.A1(_3067_),
    .A2(_3068_),
    .B1(_2913_),
    .Y(_3069_));
 sky130_fd_sc_hd__a21oi_1 _7942_ (.A1(_3066_),
    .A2(_3069_),
    .B1(_3034_),
    .Y(_3070_));
 sky130_fd_sc_hd__a221o_1 _7943_ (.A1(_2823_),
    .A2(_2853_),
    .B1(_2925_),
    .B2(net132),
    .C1(_2691_),
    .X(_3071_));
 sky130_fd_sc_hd__a221o_1 _7944_ (.A1(net106),
    .A2(_3011_),
    .B1(_3023_),
    .B2(_2763_),
    .C1(_2785_),
    .X(_3072_));
 sky130_fd_sc_hd__a31o_1 _7945_ (.A1(_2802_),
    .A2(_3071_),
    .A3(_3072_),
    .B1(_2812_),
    .X(_3073_));
 sky130_fd_sc_hd__a41o_1 _7946_ (.A1(_2923_),
    .A2(_2819_),
    .A3(_2758_),
    .A4(_2764_),
    .B1(_2679_),
    .X(_3075_));
 sky130_fd_sc_hd__o21ai_2 _7947_ (.A1(_3070_),
    .A2(_3073_),
    .B1(_3075_),
    .Y(_3076_));
 sky130_fd_sc_hd__xor2_2 _7948_ (.A(_2388_),
    .B(_2450_),
    .X(_3077_));
 sky130_fd_sc_hd__xor2_1 _7949_ (.A(_2384_),
    .B(_2452_),
    .X(_3078_));
 sky130_fd_sc_hd__mux2_1 _7950_ (.A0(_3077_),
    .A1(_3078_),
    .S(_2958_),
    .X(_3079_));
 sky130_fd_sc_hd__and3_1 _7951_ (.A(_2661_),
    .B(net118),
    .C(_3079_),
    .X(_3080_));
 sky130_fd_sc_hd__o211a_1 _7952_ (.A1(_2728_),
    .A2(_3042_),
    .B1(net113),
    .C1(_2739_),
    .X(_3081_));
 sky130_fd_sc_hd__o211a_1 _7953_ (.A1(_2728_),
    .A2(_3036_),
    .B1(net124),
    .C1(_2761_),
    .X(_3082_));
 sky130_fd_sc_hd__or3_1 _7954_ (.A(_2724_),
    .B(_3081_),
    .C(_3082_),
    .X(_3083_));
 sky130_fd_sc_hd__o21ai_1 _7955_ (.A1(_2804_),
    .A2(_2805_),
    .B1(_3045_),
    .Y(_3084_));
 sky130_fd_sc_hd__mux2_1 _7956_ (.A0(_3078_),
    .A1(_3032_),
    .S(_2958_),
    .X(_3086_));
 sky130_fd_sc_hd__mux2_1 _7957_ (.A0(_3086_),
    .A1(_3079_),
    .S(_2718_),
    .X(_3087_));
 sky130_fd_sc_hd__or4b_1 _7958_ (.A(_2769_),
    .B(_2805_),
    .C(_2728_),
    .D_N(_3087_),
    .X(_3088_));
 sky130_fd_sc_hd__a21o_1 _7959_ (.A1(_3084_),
    .A2(_3088_),
    .B1(_2918_),
    .X(_3089_));
 sky130_fd_sc_hd__a21oi_2 _7960_ (.A1(_3089_),
    .A2(_3083_),
    .B1(_3034_),
    .Y(_3090_));
 sky130_fd_sc_hd__mux4_2 _7961_ (.A0(_2915_),
    .A1(_3054_),
    .A2(_3051_),
    .A3(_3039_),
    .S0(_2855_),
    .S1(net98),
    .X(_3091_));
 sky130_fd_sc_hd__a21o_1 _7962_ (.A1(_2802_),
    .A2(_3091_),
    .B1(_2812_),
    .X(_3092_));
 sky130_fd_sc_hd__o22a_1 _7963_ (.A1(_2844_),
    .A2(_2789_),
    .B1(_3092_),
    .B2(_3090_),
    .X(_3093_));
 sky130_fd_sc_hd__a211o_1 _7964_ (.A1(_3061_),
    .A2(_3076_),
    .B1(_3093_),
    .C1(_3080_),
    .X(_3094_));
 sky130_fd_sc_hd__o211ai_2 _7965_ (.A1(_3080_),
    .A2(_3093_),
    .B1(_3061_),
    .C1(_3076_),
    .Y(_3095_));
 sky130_fd_sc_hd__and2_4 _7966_ (.A(_3094_),
    .B(_3095_),
    .X(_3097_));
 sky130_fd_sc_hd__a31o_1 _7967_ (.A1(_2923_),
    .A2(_2819_),
    .A3(_2800_),
    .B1(_2679_),
    .X(_3098_));
 sky130_fd_sc_hd__and3_1 _7968_ (.A(_2850_),
    .B(_2851_),
    .C(_2825_),
    .X(_3099_));
 sky130_fd_sc_hd__and3_1 _7969_ (.A(_2850_),
    .B(_2851_),
    .C(_2946_),
    .X(_3100_));
 sky130_fd_sc_hd__mux4_2 _7970_ (.A0(_3099_),
    .A1(_2897_),
    .A2(_3100_),
    .A3(_2941_),
    .S0(_2855_),
    .S1(net99),
    .X(_3101_));
 sky130_fd_sc_hd__a221o_1 _7971_ (.A1(_2856_),
    .A2(_2937_),
    .B1(_2939_),
    .B2(_2895_),
    .C1(_2724_),
    .X(_3102_));
 sky130_fd_sc_hd__mux2_1 _7972_ (.A0(net94),
    .A1(net93),
    .S(_2717_),
    .X(_3103_));
 sky130_fd_sc_hd__and4_1 _7973_ (.A(_2738_),
    .B(_2739_),
    .C(_2713_),
    .D(_3103_),
    .X(_3104_));
 sky130_fd_sc_hd__o211a_1 _7974_ (.A1(_2769_),
    .A2(_2771_),
    .B1(_2713_),
    .C1(_2935_),
    .X(_3105_));
 sky130_fd_sc_hd__o31a_1 _7975_ (.A1(_2786_),
    .A2(_3104_),
    .A3(_3105_),
    .B1(_2754_),
    .X(_3106_));
 sky130_fd_sc_hd__a221o_1 _7976_ (.A1(_2686_),
    .A2(_3101_),
    .B1(_3102_),
    .B2(_3106_),
    .C1(_2742_),
    .X(_3108_));
 sky130_fd_sc_hd__a22o_1 _7977_ (.A1(net93),
    .A2(_2655_),
    .B1(_3098_),
    .B2(_3108_),
    .X(_3109_));
 sky130_fd_sc_hd__nand2_1 _7978_ (.A(_2831_),
    .B(_3086_),
    .Y(_3110_));
 sky130_fd_sc_hd__or4b_1 _7979_ (.A(_2769_),
    .B(_2771_),
    .C(_2728_),
    .D_N(_2983_),
    .X(_3111_));
 sky130_fd_sc_hd__o21ai_1 _7980_ (.A1(_2804_),
    .A2(_2805_),
    .B1(_3001_),
    .Y(_3112_));
 sky130_fd_sc_hd__a21oi_2 _7981_ (.A1(_3111_),
    .A2(_3112_),
    .B1(_2786_),
    .Y(_3113_));
 sky130_fd_sc_hd__o21a_1 _7982_ (.A1(_2881_),
    .A2(_2890_),
    .B1(_2786_),
    .X(_3114_));
 sky130_fd_sc_hd__a21o_1 _7983_ (.A1(net113),
    .A2(_2739_),
    .B1(_2972_),
    .X(_3115_));
 sky130_fd_sc_hd__mux2_1 _7984_ (.A0(_3033_),
    .A1(_3086_),
    .S(_2718_),
    .X(_3116_));
 sky130_fd_sc_hd__or4b_1 _7985_ (.A(_2804_),
    .B(_2805_),
    .C(_2728_),
    .D_N(_3116_),
    .X(_3117_));
 sky130_fd_sc_hd__a21oi_1 _7986_ (.A1(_3115_),
    .A2(_3117_),
    .B1(_2918_),
    .Y(_3119_));
 sky130_fd_sc_hd__a22o_1 _7987_ (.A1(net123),
    .A2(_2761_),
    .B1(_3014_),
    .B2(_2963_),
    .X(_3120_));
 sky130_fd_sc_hd__a2bb2o_1 _7988_ (.A1_N(_2728_),
    .A2_N(_2993_),
    .B1(_2738_),
    .B2(_2739_),
    .X(_3121_));
 sky130_fd_sc_hd__a31o_1 _7989_ (.A1(_2880_),
    .A2(_3120_),
    .A3(_3121_),
    .B1(_2686_),
    .X(_3122_));
 sky130_fd_sc_hd__o32a_1 _7990_ (.A1(_2756_),
    .A2(_3113_),
    .A3(_3114_),
    .B1(_3119_),
    .B2(_3122_),
    .X(_3123_));
 sky130_fd_sc_hd__o2bb2ai_2 _7991_ (.A1_N(_2746_),
    .A2_N(_2811_),
    .B1(_3123_),
    .B2(_2812_),
    .Y(_3124_));
 sky130_fd_sc_hd__nand3_2 _7992_ (.A(_3109_),
    .B(_3110_),
    .C(_3124_),
    .Y(_3125_));
 sky130_fd_sc_hd__a21o_1 _7993_ (.A1(_3110_),
    .A2(_3124_),
    .B1(_3109_),
    .X(_3126_));
 sky130_fd_sc_hd__and2_1 _7994_ (.A(_3125_),
    .B(_3126_),
    .X(_3127_));
 sky130_fd_sc_hd__nand4_2 _7995_ (.A(_3010_),
    .B(_3060_),
    .C(_3097_),
    .D(_3127_),
    .Y(_3128_));
 sky130_fd_sc_hd__o21ai_1 _7996_ (.A1(_3027_),
    .A2(_2827_),
    .B1(_2820_),
    .Y(_3130_));
 sky130_fd_sc_hd__a221o_1 _7997_ (.A1(_2824_),
    .A2(_2897_),
    .B1(_2946_),
    .B2(_2716_),
    .C1(_2724_),
    .X(_3131_));
 sky130_fd_sc_hd__a221o_1 _7998_ (.A1(_2939_),
    .A2(_2716_),
    .B1(_2941_),
    .B2(_2823_),
    .C1(_2786_),
    .X(_3132_));
 sky130_fd_sc_hd__a221o_1 _7999_ (.A1(_2917_),
    .A2(_2935_),
    .B1(_2937_),
    .B2(_2824_),
    .C1(_2803_),
    .X(_3133_));
 sky130_fd_sc_hd__mux2_1 _8000_ (.A0(net92),
    .A1(net91),
    .S(_2729_),
    .X(_3134_));
 sky130_fd_sc_hd__and3_1 _8001_ (.A(_2850_),
    .B(_2851_),
    .C(_3134_),
    .X(_3135_));
 sky130_fd_sc_hd__a221o_1 _8002_ (.A1(_2895_),
    .A2(_3103_),
    .B1(_3135_),
    .B2(_2856_),
    .C1(_2918_),
    .X(_3136_));
 sky130_fd_sc_hd__a31o_1 _8003_ (.A1(_2923_),
    .A2(_3133_),
    .A3(_3136_),
    .B1(_2812_),
    .X(_3137_));
 sky130_fd_sc_hd__a31o_1 _8004_ (.A1(_2687_),
    .A2(_3131_),
    .A3(_3132_),
    .B1(_3137_),
    .X(_3138_));
 sky130_fd_sc_hd__a22o_1 _8005_ (.A1(net91),
    .A2(_2658_),
    .B1(_3130_),
    .B2(_3138_),
    .X(_3139_));
 sky130_fd_sc_hd__xor2_2 _8006_ (.A(_2393_),
    .B(_2448_),
    .X(_3141_));
 sky130_fd_sc_hd__mux2_1 _8007_ (.A0(_3141_),
    .A1(_3077_),
    .S(_2958_),
    .X(_3142_));
 sky130_fd_sc_hd__mux2_1 _8008_ (.A0(_3079_),
    .A1(_3142_),
    .S(_2794_),
    .X(_3143_));
 sky130_fd_sc_hd__and2_1 _8009_ (.A(_2917_),
    .B(_3143_),
    .X(_3144_));
 sky130_fd_sc_hd__a31o_1 _8010_ (.A1(_2824_),
    .A2(_3014_),
    .A3(_3116_),
    .B1(_2913_),
    .X(_3145_));
 sky130_fd_sc_hd__o2bb2a_1 _8011_ (.A1_N(_2913_),
    .A2_N(_2973_),
    .B1(_3144_),
    .B2(_3145_),
    .X(_3146_));
 sky130_fd_sc_hd__nor2_1 _8012_ (.A(_2687_),
    .B(_3146_),
    .Y(_3147_));
 sky130_fd_sc_hd__nand3_1 _8013_ (.A(_2918_),
    .B(_3002_),
    .C(_3003_),
    .Y(_3148_));
 sky130_fd_sc_hd__o211a_1 _8014_ (.A1(_2913_),
    .A2(_2995_),
    .B1(_3148_),
    .C1(_2687_),
    .X(_3149_));
 sky130_fd_sc_hd__and3_1 _8015_ (.A(net130),
    .B(_2742_),
    .C(_2676_),
    .X(_3150_));
 sky130_fd_sc_hd__a22oi_1 _8016_ (.A1(_2831_),
    .A2(_3142_),
    .B1(_3150_),
    .B2(_2841_),
    .Y(_3152_));
 sky130_fd_sc_hd__o31a_2 _8017_ (.A1(_2746_),
    .A2(_3147_),
    .A3(_3149_),
    .B1(_3152_),
    .X(_3153_));
 sky130_fd_sc_hd__nor2_1 _8018_ (.A(_3139_),
    .B(_3153_),
    .Y(_3154_));
 sky130_fd_sc_hd__a31o_1 _8019_ (.A1(_2923_),
    .A2(_2894_),
    .A3(_2899_),
    .B1(_2670_),
    .X(_3155_));
 sky130_fd_sc_hd__and3_1 _8020_ (.A(_2850_),
    .B(_2851_),
    .C(_2939_),
    .X(_3156_));
 sky130_fd_sc_hd__mux4_2 _8021_ (.A0(_3100_),
    .A1(_3156_),
    .A2(_2941_),
    .A3(_2937_),
    .S0(_2692_),
    .S1(_2856_),
    .X(_3157_));
 sky130_fd_sc_hd__or3_4 _8022_ (.A(_2692_),
    .B(_3104_),
    .C(_3105_),
    .X(_3158_));
 sky130_fd_sc_hd__mux2_1 _8023_ (.A0(net88),
    .A1(net77),
    .S(_2730_),
    .X(_3159_));
 sky130_fd_sc_hd__and4_1 _8024_ (.A(_2738_),
    .B(_2739_),
    .C(_2713_),
    .D(_3159_),
    .X(_3160_));
 sky130_fd_sc_hd__and3_1 _8025_ (.A(_2760_),
    .B(_2761_),
    .C(_3135_),
    .X(_3161_));
 sky130_fd_sc_hd__o31a_1 _8026_ (.A1(_2786_),
    .A2(_3160_),
    .A3(_3161_),
    .B1(_2754_),
    .X(_3163_));
 sky130_fd_sc_hd__a221o_1 _8027_ (.A1(_3157_),
    .A2(_2802_),
    .B1(_3158_),
    .B2(_3163_),
    .C1(_2742_),
    .X(_3164_));
 sky130_fd_sc_hd__a32o_2 _8028_ (.A1(_3164_),
    .A2(_3155_),
    .A3(_2819_),
    .B1(_2657_),
    .B2(net77),
    .X(_3165_));
 sky130_fd_sc_hd__nand3_1 _8029_ (.A(_2913_),
    .B(_3111_),
    .C(_3112_),
    .Y(_3166_));
 sky130_fd_sc_hd__a21o_1 _8030_ (.A1(_3120_),
    .A2(_3121_),
    .B1(_2918_),
    .X(_3167_));
 sky130_fd_sc_hd__nand3_1 _8031_ (.A(_2913_),
    .B(_3115_),
    .C(_3117_),
    .Y(_3168_));
 sky130_fd_sc_hd__o211a_1 _8032_ (.A1(_2804_),
    .A2(_2805_),
    .B1(_3014_),
    .C1(_3143_),
    .X(_3169_));
 sky130_fd_sc_hd__or2b_1 _8033_ (.A(_2446_),
    .B_N(_2398_),
    .X(_3170_));
 sky130_fd_sc_hd__xnor2_2 _8034_ (.A(_3170_),
    .B(_2445_),
    .Y(_3171_));
 sky130_fd_sc_hd__mux2_1 _8035_ (.A0(_3171_),
    .A1(_3141_),
    .S(_2958_),
    .X(_3172_));
 sky130_fd_sc_hd__xor2_2 _8036_ (.A(_2439_),
    .B(_2443_),
    .X(_3174_));
 sky130_fd_sc_hd__mux2_1 _8037_ (.A0(_3174_),
    .A1(_3171_),
    .S(_2958_),
    .X(_3175_));
 sky130_fd_sc_hd__mux2_1 _8038_ (.A0(_3172_),
    .A1(_3175_),
    .S(_2794_),
    .X(_3176_));
 sky130_fd_sc_hd__and4_1 _8039_ (.A(net113),
    .B(_2739_),
    .C(_3014_),
    .D(_3176_),
    .X(_3177_));
 sky130_fd_sc_hd__o31a_1 _8040_ (.A1(_2880_),
    .A2(_3169_),
    .A3(_3177_),
    .B1(_2756_),
    .X(_3178_));
 sky130_fd_sc_hd__a32o_1 _8041_ (.A1(_3034_),
    .A2(_3166_),
    .A3(_3167_),
    .B1(_3168_),
    .B2(_3178_),
    .X(_3179_));
 sky130_fd_sc_hd__and3_1 _8042_ (.A(_2661_),
    .B(net118),
    .C(_3175_),
    .X(_3180_));
 sky130_fd_sc_hd__a41o_1 _8043_ (.A1(_2923_),
    .A2(_2879_),
    .A3(_2891_),
    .A4(_3150_),
    .B1(_3180_),
    .X(_3181_));
 sky130_fd_sc_hd__a21oi_4 _8044_ (.A1(_2844_),
    .A2(_3179_),
    .B1(_3181_),
    .Y(_3182_));
 sky130_fd_sc_hd__or2_4 _8045_ (.A(_3165_),
    .B(_3182_),
    .X(_3183_));
 sky130_fd_sc_hd__and2_1 _8046_ (.A(net66),
    .B(_2657_),
    .X(_3185_));
 sky130_fd_sc_hd__a221o_1 _8047_ (.A1(_2917_),
    .A2(_3011_),
    .B1(_3023_),
    .B2(_2895_),
    .C1(_2803_),
    .X(_3186_));
 sky130_fd_sc_hd__or3_1 _8048_ (.A(_2880_),
    .B(_3067_),
    .C(_3068_),
    .X(_3187_));
 sky130_fd_sc_hd__and3_1 _8049_ (.A(_3034_),
    .B(_3186_),
    .C(_3187_),
    .X(_3188_));
 sky130_fd_sc_hd__or3_1 _8050_ (.A(_2803_),
    .B(_3062_),
    .C(_3065_),
    .X(_3189_));
 sky130_fd_sc_hd__mux2_1 _8051_ (.A0(net91),
    .A1(net88),
    .S(_2718_),
    .X(_3190_));
 sky130_fd_sc_hd__and3_1 _8052_ (.A(_2850_),
    .B(_2851_),
    .C(_3190_),
    .X(_3191_));
 sky130_fd_sc_hd__mux2_1 _8053_ (.A0(net77),
    .A1(net66),
    .S(_2794_),
    .X(_3192_));
 sky130_fd_sc_hd__a221o_1 _8054_ (.A1(_2824_),
    .A2(_3191_),
    .B1(_3192_),
    .B2(_2917_),
    .C1(_2918_),
    .X(_3193_));
 sky130_fd_sc_hd__a31o_1 _8055_ (.A1(_2835_),
    .A2(_3189_),
    .A3(_3193_),
    .B1(_2812_),
    .X(_3194_));
 sky130_fd_sc_hd__o22a_2 _8056_ (.A1(_2680_),
    .A2(_2927_),
    .B1(_3188_),
    .B2(_3194_),
    .X(_3196_));
 sky130_fd_sc_hd__a221o_1 _8057_ (.A1(_2895_),
    .A2(_3050_),
    .B1(_3039_),
    .B2(_2856_),
    .C1(_2758_),
    .X(_3197_));
 sky130_fd_sc_hd__o21ai_1 _8058_ (.A1(_3081_),
    .A2(_3082_),
    .B1(_2758_),
    .Y(_3198_));
 sky130_fd_sc_hd__a21o_1 _8059_ (.A1(_3197_),
    .A2(_3198_),
    .B1(_2757_),
    .X(_3199_));
 sky130_fd_sc_hd__mux2_1 _8060_ (.A0(_3142_),
    .A1(_3172_),
    .S(_2794_),
    .X(_3200_));
 sky130_fd_sc_hd__xor2_2 _8061_ (.A(_2402_),
    .B(_2437_),
    .X(_3201_));
 sky130_fd_sc_hd__mux2_1 _8062_ (.A0(_3201_),
    .A1(_3174_),
    .S(_2958_),
    .X(_3202_));
 sky130_fd_sc_hd__mux2_1 _8063_ (.A0(_3175_),
    .A1(_3202_),
    .S(_2794_),
    .X(_3203_));
 sky130_fd_sc_hd__a22o_1 _8064_ (.A1(_2895_),
    .A2(_3200_),
    .B1(_3203_),
    .B2(_2917_),
    .X(_3204_));
 sky130_fd_sc_hd__a21oi_1 _8065_ (.A1(_3084_),
    .A2(_3088_),
    .B1(_2758_),
    .Y(_3205_));
 sky130_fd_sc_hd__a211o_1 _8066_ (.A1(_2758_),
    .A2(_3204_),
    .B1(_3205_),
    .C1(_2687_),
    .X(_3207_));
 sky130_fd_sc_hd__and3_1 _8067_ (.A(_2661_),
    .B(net118),
    .C(_3202_),
    .X(_3208_));
 sky130_fd_sc_hd__a41o_1 _8068_ (.A1(_2757_),
    .A2(_2914_),
    .A3(_2919_),
    .A4(_3150_),
    .B1(_3208_),
    .X(_3209_));
 sky130_fd_sc_hd__a31oi_4 _8069_ (.A1(_2844_),
    .A2(_3199_),
    .A3(_3207_),
    .B1(_3209_),
    .Y(_3210_));
 sky130_fd_sc_hd__a2111o_1 _8070_ (.A1(_3182_),
    .A2(_3165_),
    .B1(_3185_),
    .C1(_3196_),
    .D1(_3210_),
    .X(_3211_));
 sky130_fd_sc_hd__nand2_1 _8071_ (.A(net88),
    .B(_2658_),
    .Y(_3212_));
 sky130_fd_sc_hd__a221o_1 _8072_ (.A1(_2895_),
    .A2(_2925_),
    .B1(_3023_),
    .B2(net132),
    .C1(net100),
    .X(_3213_));
 sky130_fd_sc_hd__a221o_1 _8073_ (.A1(_2763_),
    .A2(_3011_),
    .B1(_3012_),
    .B2(net132),
    .C1(_2786_),
    .X(_3214_));
 sky130_fd_sc_hd__and3_1 _8074_ (.A(_3034_),
    .B(_3213_),
    .C(_3214_),
    .X(_3215_));
 sky130_fd_sc_hd__a221o_1 _8075_ (.A1(_2895_),
    .A2(_3064_),
    .B1(_3191_),
    .B2(_2856_),
    .C1(_2918_),
    .X(_3216_));
 sky130_fd_sc_hd__o311a_1 _8076_ (.A1(_2758_),
    .A2(_3016_),
    .A3(_3018_),
    .B1(_3216_),
    .C1(_2835_),
    .X(_3218_));
 sky130_fd_sc_hd__a41o_1 _8077_ (.A1(_2757_),
    .A2(_2819_),
    .A3(_2849_),
    .A4(_2857_),
    .B1(_2680_),
    .X(_3219_));
 sky130_fd_sc_hd__o31ai_4 _8078_ (.A1(_2812_),
    .A2(_3215_),
    .A3(_3218_),
    .B1(_3219_),
    .Y(_3220_));
 sky130_fd_sc_hd__and2_1 _8079_ (.A(_3014_),
    .B(_3087_),
    .X(_3221_));
 sky130_fd_sc_hd__a22o_1 _8080_ (.A1(_2824_),
    .A2(_3221_),
    .B1(_3200_),
    .B2(_2917_),
    .X(_3222_));
 sky130_fd_sc_hd__o211a_1 _8081_ (.A1(_2856_),
    .A2(_3043_),
    .B1(_3046_),
    .C1(_2918_),
    .X(_3223_));
 sky130_fd_sc_hd__a211o_1 _8082_ (.A1(_2758_),
    .A2(_3222_),
    .B1(_3223_),
    .C1(_3034_),
    .X(_3224_));
 sky130_fd_sc_hd__a21o_1 _8083_ (.A1(_3053_),
    .A2(_3055_),
    .B1(_2803_),
    .X(_3225_));
 sky130_fd_sc_hd__a221o_1 _8084_ (.A1(_2716_),
    .A2(_3037_),
    .B1(_3039_),
    .B2(_2824_),
    .C1(_2880_),
    .X(_3226_));
 sky130_fd_sc_hd__a21o_1 _8085_ (.A1(_3225_),
    .A2(_3226_),
    .B1(_2835_),
    .X(_3227_));
 sky130_fd_sc_hd__and3_1 _8086_ (.A(_2661_),
    .B(net118),
    .C(_3172_),
    .X(_3229_));
 sky130_fd_sc_hd__a41o_1 _8087_ (.A1(_2835_),
    .A2(_2860_),
    .A3(_2871_),
    .A4(_3150_),
    .B1(_3229_),
    .X(_3230_));
 sky130_fd_sc_hd__a31o_1 _8088_ (.A1(_2844_),
    .A2(_3224_),
    .A3(_3227_),
    .B1(_3230_),
    .X(_3231_));
 sky130_fd_sc_hd__nand3_1 _8089_ (.A(_3212_),
    .B(_3220_),
    .C(_3231_),
    .Y(_3232_));
 sky130_fd_sc_hd__a21oi_4 _8090_ (.A1(_3212_),
    .A2(_3220_),
    .B1(_3231_),
    .Y(_3233_));
 sky130_fd_sc_hd__a31oi_2 _8091_ (.A1(_3211_),
    .A2(_3183_),
    .A3(_3232_),
    .B1(_3233_),
    .Y(_3234_));
 sky130_fd_sc_hd__nand2_1 _8092_ (.A(_3139_),
    .B(_3153_),
    .Y(_3235_));
 sky130_fd_sc_hd__o21a_1 _8093_ (.A1(_3234_),
    .A2(_3154_),
    .B1(_3235_),
    .X(_3236_));
 sky130_fd_sc_hd__and2_1 _8094_ (.A(_2954_),
    .B(_3009_),
    .X(_3237_));
 sky130_fd_sc_hd__a21bo_1 _8095_ (.A1(_3125_),
    .A2(_3094_),
    .B1_N(_3126_),
    .X(_3238_));
 sky130_fd_sc_hd__or2_1 _8096_ (.A(_2954_),
    .B(_3009_),
    .X(_3240_));
 sky130_fd_sc_hd__nand4bb_1 _8097_ (.A_N(_3237_),
    .B_N(_3238_),
    .C(_3240_),
    .D(_3060_),
    .Y(_3241_));
 sky130_fd_sc_hd__a22o_1 _8098_ (.A1(net94),
    .A2(_2658_),
    .B1(_3026_),
    .B2(_3028_),
    .X(_3242_));
 sky130_fd_sc_hd__and2_1 _8099_ (.A(_3242_),
    .B(_3059_),
    .X(_3243_));
 sky130_fd_sc_hd__o21ai_1 _8100_ (.A1(_3237_),
    .A2(_3243_),
    .B1(_3240_),
    .Y(_3244_));
 sky130_fd_sc_hd__o211ai_2 _8101_ (.A1(_3236_),
    .A2(_3128_),
    .B1(_3241_),
    .C1(_3244_),
    .Y(_3245_));
 sky130_fd_sc_hd__a21o_1 _8102_ (.A1(_3186_),
    .A2(_3187_),
    .B1(_3034_),
    .X(_3246_));
 sky130_fd_sc_hd__a21o_1 _8103_ (.A1(_2924_),
    .A2(_2926_),
    .B1(_2835_),
    .X(_3247_));
 sky130_fd_sc_hd__a32o_1 _8104_ (.A1(_2680_),
    .A2(_3246_),
    .A3(_3247_),
    .B1(_2657_),
    .B2(net96),
    .X(_3248_));
 sky130_fd_sc_hd__a21oi_1 _8105_ (.A1(_2914_),
    .A2(_2919_),
    .B1(_2835_),
    .Y(_3249_));
 sky130_fd_sc_hd__a21oi_1 _8106_ (.A1(_3197_),
    .A2(_3198_),
    .B1(_2687_),
    .Y(_3251_));
 sky130_fd_sc_hd__o32a_1 _8107_ (.A1(_2746_),
    .A2(_3249_),
    .A3(_3251_),
    .B1(_2967_),
    .B2(_2747_),
    .X(_3252_));
 sky130_fd_sc_hd__nand2_1 _8108_ (.A(_3248_),
    .B(_3252_),
    .Y(_3253_));
 sky130_fd_sc_hd__or2_1 _8109_ (.A(_3248_),
    .B(_3252_),
    .X(_3254_));
 sky130_fd_sc_hd__nand2_2 _8110_ (.A(_3253_),
    .B(_3254_),
    .Y(_3255_));
 sky130_fd_sc_hd__or2_1 _8111_ (.A(_2802_),
    .B(_3157_),
    .X(_3256_));
 sky130_fd_sc_hd__a21o_1 _8112_ (.A1(_2894_),
    .A2(_2899_),
    .B1(_2923_),
    .X(_3257_));
 sky130_fd_sc_hd__a32o_2 _8113_ (.A1(_2680_),
    .A2(_3256_),
    .A3(_3257_),
    .B1(_2657_),
    .B2(net97),
    .X(_3258_));
 sky130_fd_sc_hd__a21oi_1 _8114_ (.A1(_3166_),
    .A2(_3167_),
    .B1(_3034_),
    .Y(_3259_));
 sky130_fd_sc_hd__a21oi_1 _8115_ (.A1(_2879_),
    .A2(_2891_),
    .B1(_2835_),
    .Y(_3260_));
 sky130_fd_sc_hd__o32a_1 _8116_ (.A1(_2746_),
    .A2(_3259_),
    .A3(_3260_),
    .B1(_2961_),
    .B2(_2747_),
    .X(_3262_));
 sky130_fd_sc_hd__nand2_1 _8117_ (.A(_3258_),
    .B(_3262_),
    .Y(_3263_));
 sky130_fd_sc_hd__or2_1 _8118_ (.A(_3258_),
    .B(_3262_),
    .X(_3264_));
 sky130_fd_sc_hd__nand2_4 _8119_ (.A(_3263_),
    .B(_3264_),
    .Y(_3265_));
 sky130_fd_sc_hd__nor2_1 _8120_ (.A(_3255_),
    .B(_3265_),
    .Y(_3266_));
 sky130_fd_sc_hd__a21o_1 _8121_ (.A1(_2945_),
    .A2(_2947_),
    .B1(_2686_),
    .X(_3267_));
 sky130_fd_sc_hd__a31o_1 _8122_ (.A1(_2794_),
    .A2(_2724_),
    .A3(_2716_),
    .B1(_2754_),
    .X(_3268_));
 sky130_fd_sc_hd__a32o_2 _8123_ (.A1(_2679_),
    .A2(_3267_),
    .A3(_3268_),
    .B1(_2655_),
    .B2(net72),
    .X(_3269_));
 sky130_fd_sc_hd__o21ai_1 _8124_ (.A1(_2998_),
    .A2(_3004_),
    .B1(_2756_),
    .Y(_3270_));
 sky130_fd_sc_hd__a32o_2 _8125_ (.A1(_3270_),
    .A2(_3268_),
    .A3(_2844_),
    .B1(_2999_),
    .B2(_2830_),
    .X(_3271_));
 sky130_fd_sc_hd__xor2_4 _8126_ (.A(_3271_),
    .B(_3269_),
    .X(_3273_));
 sky130_fd_sc_hd__a21o_1 _8127_ (.A1(_3022_),
    .A2(_3024_),
    .B1(_2685_),
    .X(_3274_));
 sky130_fd_sc_hd__nand2_1 _8128_ (.A(_2686_),
    .B(_2720_),
    .Y(_3275_));
 sky130_fd_sc_hd__a32o_4 _8129_ (.A1(_2679_),
    .A2(_3274_),
    .A3(_3275_),
    .B1(_2655_),
    .B2(net71),
    .X(_3276_));
 sky130_fd_sc_hd__a21o_1 _8130_ (.A1(_3049_),
    .A2(_3056_),
    .B1(_2686_),
    .X(_3277_));
 sky130_fd_sc_hd__nand2_1 _8131_ (.A(_2686_),
    .B(_2741_),
    .Y(_3278_));
 sky130_fd_sc_hd__a32oi_4 _8132_ (.A1(_3278_),
    .A2(_3277_),
    .A3(_2842_),
    .B1(_2977_),
    .B2(_2830_),
    .Y(_3279_));
 sky130_fd_sc_hd__xnor2_4 _8133_ (.A(_3279_),
    .B(_3276_),
    .Y(_3280_));
 sky130_fd_sc_hd__a21o_1 _8134_ (.A1(_3071_),
    .A2(_3072_),
    .B1(_2685_),
    .X(_3281_));
 sky130_fd_sc_hd__a21o_1 _8135_ (.A1(_2724_),
    .A2(_2764_),
    .B1(_2754_),
    .X(_3282_));
 sky130_fd_sc_hd__a32o_4 _8136_ (.A1(_2679_),
    .A2(_3281_),
    .A3(_3282_),
    .B1(_2655_),
    .B2(net69),
    .X(_3284_));
 sky130_fd_sc_hd__mux2_1 _8137_ (.A0(_2787_),
    .A1(_3091_),
    .S(_2754_),
    .X(_3285_));
 sky130_fd_sc_hd__o2bb2a_2 _8138_ (.A1_N(_2844_),
    .A2_N(_3285_),
    .B1(_2990_),
    .B2(_2747_),
    .X(_3286_));
 sky130_fd_sc_hd__xor2_4 _8139_ (.A(_3286_),
    .B(_3284_),
    .X(_3287_));
 sky130_fd_sc_hd__mux2_1 _8140_ (.A0(_2800_),
    .A1(_3101_),
    .S(_2754_),
    .X(_3288_));
 sky130_fd_sc_hd__a22o_4 _8141_ (.A1(net70),
    .A2(_2655_),
    .B1(_2679_),
    .B2(_3288_),
    .X(_3289_));
 sky130_fd_sc_hd__nand2_1 _8142_ (.A(_2802_),
    .B(_2809_),
    .Y(_3290_));
 sky130_fd_sc_hd__o31a_1 _8143_ (.A1(_2686_),
    .A2(_3113_),
    .A3(_3114_),
    .B1(_2842_),
    .X(_3291_));
 sky130_fd_sc_hd__o2bb2a_4 _8144_ (.A1_N(_3290_),
    .A2_N(_3291_),
    .B1(_2747_),
    .B2(_2981_),
    .X(_3292_));
 sky130_fd_sc_hd__xor2_4 _8145_ (.A(_3289_),
    .B(_3292_),
    .X(_3293_));
 sky130_fd_sc_hd__nand4bb_4 _8146_ (.A_N(_3273_),
    .B_N(_3280_),
    .C(_3287_),
    .D(_3293_),
    .Y(_3295_));
 sky130_fd_sc_hd__inv_2 _8147_ (.A(_3295_),
    .Y(_3296_));
 sky130_fd_sc_hd__a21o_1 _8148_ (.A1(_3131_),
    .A2(_3132_),
    .B1(_2802_),
    .X(_3297_));
 sky130_fd_sc_hd__a21o_1 _8149_ (.A1(_2822_),
    .A2(_2826_),
    .B1(_2756_),
    .X(_3298_));
 sky130_fd_sc_hd__a32o_2 _8150_ (.A1(_3297_),
    .A2(_2680_),
    .A3(_3298_),
    .B1(_2657_),
    .B2(net68),
    .X(_3299_));
 sky130_fd_sc_hd__o211a_1 _8151_ (.A1(_2913_),
    .A2(_2995_),
    .B1(_3148_),
    .C1(_2756_),
    .X(_3300_));
 sky130_fd_sc_hd__a21oi_1 _8152_ (.A1(_2822_),
    .A2(_2840_),
    .B1(_2923_),
    .Y(_3301_));
 sky130_fd_sc_hd__o32a_2 _8153_ (.A1(_2746_),
    .A2(_3300_),
    .A3(_3301_),
    .B1(_2992_),
    .B2(_2747_),
    .X(_3302_));
 sky130_fd_sc_hd__xnor2_4 _8154_ (.A(_3302_),
    .B(_3299_),
    .Y(_3303_));
 sky130_fd_sc_hd__a21o_1 _8155_ (.A1(_3213_),
    .A2(_3214_),
    .B1(_2802_),
    .X(_3304_));
 sky130_fd_sc_hd__a21o_1 _8156_ (.A1(_2849_),
    .A2(_2857_),
    .B1(_2756_),
    .X(_3306_));
 sky130_fd_sc_hd__a32o_4 _8157_ (.A1(_2679_),
    .A2(_3304_),
    .A3(_3306_),
    .B1(_2655_),
    .B2(net67),
    .X(_3307_));
 sky130_fd_sc_hd__a21oi_1 _8158_ (.A1(_2860_),
    .A2(_2871_),
    .B1(_2923_),
    .Y(_3308_));
 sky130_fd_sc_hd__a21oi_1 _8159_ (.A1(_3225_),
    .A2(_3226_),
    .B1(_3034_),
    .Y(_3309_));
 sky130_fd_sc_hd__o32a_4 _8160_ (.A1(_2746_),
    .A2(_3308_),
    .A3(_3309_),
    .B1(_2959_),
    .B2(_2747_),
    .X(_3310_));
 sky130_fd_sc_hd__xnor2_4 _8161_ (.A(_3307_),
    .B(_3310_),
    .Y(_3311_));
 sky130_fd_sc_hd__nor2_1 _8162_ (.A(_3303_),
    .B(_3311_),
    .Y(_3312_));
 sky130_fd_sc_hd__and3_1 _8163_ (.A(_3266_),
    .B(_3296_),
    .C(_3312_),
    .X(_3313_));
 sky130_fd_sc_hd__nand2_1 _8164_ (.A(_3299_),
    .B(_3302_),
    .Y(_3314_));
 sky130_fd_sc_hd__nand2_1 _8165_ (.A(_3307_),
    .B(_3310_),
    .Y(_3315_));
 sky130_fd_sc_hd__nor2_1 _8166_ (.A(_3299_),
    .B(_3302_),
    .Y(_3317_));
 sky130_fd_sc_hd__a21o_1 _8167_ (.A1(_3314_),
    .A2(_3315_),
    .B1(_3317_),
    .X(_3318_));
 sky130_fd_sc_hd__nor2_1 _8168_ (.A(_3273_),
    .B(_3280_),
    .Y(_3319_));
 sky130_fd_sc_hd__nand2_1 _8169_ (.A(_3284_),
    .B(_3286_),
    .Y(_3320_));
 sky130_fd_sc_hd__nand2_1 _8170_ (.A(_3289_),
    .B(_3292_),
    .Y(_3321_));
 sky130_fd_sc_hd__nor2_1 _8171_ (.A(_3289_),
    .B(_3292_),
    .Y(_3322_));
 sky130_fd_sc_hd__a21oi_1 _8172_ (.A1(_3320_),
    .A2(_3321_),
    .B1(_3322_),
    .Y(_3323_));
 sky130_fd_sc_hd__nand2b_1 _8173_ (.A_N(_3269_),
    .B(_3271_),
    .Y(_3324_));
 sky130_fd_sc_hd__and3_1 _8174_ (.A(_3324_),
    .B(_3276_),
    .C(_3279_),
    .X(_3325_));
 sky130_fd_sc_hd__and2b_1 _8175_ (.A_N(_3271_),
    .B(_3269_),
    .X(_3326_));
 sky130_fd_sc_hd__a211oi_1 _8176_ (.A1(_3319_),
    .A2(_3323_),
    .B1(_3325_),
    .C1(_3326_),
    .Y(_3328_));
 sky130_fd_sc_hd__or2_4 _8177_ (.A(_3303_),
    .B(_3311_),
    .X(_3329_));
 sky130_fd_sc_hd__a21bo_1 _8178_ (.A1(_3253_),
    .A2(_3263_),
    .B1_N(_3264_),
    .X(_3330_));
 sky130_fd_sc_hd__or3_4 _8179_ (.A(_3295_),
    .B(_3329_),
    .C(_3330_),
    .X(_3331_));
 sky130_fd_sc_hd__o211ai_2 _8180_ (.A1(_3295_),
    .A2(_3318_),
    .B1(_3328_),
    .C1(_3331_),
    .Y(_3332_));
 sky130_fd_sc_hd__a21o_1 _8181_ (.A1(_3313_),
    .A2(_3245_),
    .B1(_3332_),
    .X(_3333_));
 sky130_fd_sc_hd__nand2_1 _8182_ (.A(_2846_),
    .B(_2874_),
    .Y(_3334_));
 sky130_fd_sc_hd__inv_2 _8183_ (.A(_2929_),
    .Y(_3335_));
 sky130_fd_sc_hd__o21a_1 _8184_ (.A1(_2902_),
    .A2(_3335_),
    .B1(_2903_),
    .X(_3336_));
 sky130_fd_sc_hd__a22o_1 _8185_ (.A1(_2847_),
    .A2(_3334_),
    .B1(_2878_),
    .B2(_3336_),
    .X(_3337_));
 sky130_fd_sc_hd__a21oi_4 _8186_ (.A1(_3333_),
    .A2(_2934_),
    .B1(_3337_),
    .Y(_3339_));
 sky130_fd_sc_hd__a21o_1 _8187_ (.A1(_2791_),
    .A2(_2815_),
    .B1(_2814_),
    .X(_3340_));
 sky130_fd_sc_hd__and3_1 _8188_ (.A(_2748_),
    .B(_2723_),
    .C(_2749_),
    .X(_3341_));
 sky130_fd_sc_hd__or2_1 _8189_ (.A(_2658_),
    .B(_3341_),
    .X(_3342_));
 sky130_fd_sc_hd__o21ba_2 _8190_ (.A1(_2753_),
    .A2(_3340_),
    .B1_N(_3342_),
    .X(_3343_));
 sky130_fd_sc_hd__o21a_4 _8191_ (.A1(_3339_),
    .A2(_2818_),
    .B1(_3343_),
    .X(_3344_));
 sky130_fd_sc_hd__buf_4 _8192_ (.A(_3344_),
    .X(_3345_));
 sky130_fd_sc_hd__xnor2_2 _8193_ (.A(\In2_reg[31] ),
    .B(\In1_reg[31] ),
    .Y(_3346_));
 sky130_fd_sc_hd__nand2_1 _8194_ (.A(_3345_),
    .B(_3346_),
    .Y(_3347_));
 sky130_fd_sc_hd__buf_2 _8195_ (.A(net65),
    .X(_3348_));
 sky130_fd_sc_hd__buf_2 _8196_ (.A(_3348_),
    .X(_3350_));
 sky130_fd_sc_hd__o211a_1 _8197_ (.A1(\F1.sign_b ),
    .A2(_3345_),
    .B1(_3347_),
    .C1(_3350_),
    .X(_0032_));
 sky130_fd_sc_hd__and2_1 _8198_ (.A(_2276_),
    .B(net33),
    .X(_3351_));
 sky130_fd_sc_hd__clkbuf_1 _8199_ (.A(_3351_),
    .X(_0033_));
 sky130_fd_sc_hd__and2_1 _8200_ (.A(_2276_),
    .B(net44),
    .X(_3352_));
 sky130_fd_sc_hd__clkbuf_1 _8201_ (.A(_3352_),
    .X(_0034_));
 sky130_fd_sc_hd__and2_1 _8202_ (.A(_2276_),
    .B(net55),
    .X(_3353_));
 sky130_fd_sc_hd__clkbuf_1 _8203_ (.A(_3353_),
    .X(_0035_));
 sky130_fd_sc_hd__and2_1 _8204_ (.A(_2276_),
    .B(net58),
    .X(_3354_));
 sky130_fd_sc_hd__clkbuf_1 _8205_ (.A(_3354_),
    .X(_0036_));
 sky130_fd_sc_hd__and2_1 _8206_ (.A(_2276_),
    .B(net59),
    .X(_3356_));
 sky130_fd_sc_hd__clkbuf_1 _8207_ (.A(_3356_),
    .X(_0037_));
 sky130_fd_sc_hd__clkbuf_2 _8208_ (.A(net65),
    .X(_3357_));
 sky130_fd_sc_hd__and2_1 _8209_ (.A(_3357_),
    .B(net60),
    .X(_3358_));
 sky130_fd_sc_hd__clkbuf_1 _8210_ (.A(_3358_),
    .X(_0038_));
 sky130_fd_sc_hd__and2_1 _8211_ (.A(_3357_),
    .B(net61),
    .X(_3359_));
 sky130_fd_sc_hd__clkbuf_1 _8212_ (.A(_3359_),
    .X(_0039_));
 sky130_fd_sc_hd__and2_1 _8213_ (.A(_3357_),
    .B(net62),
    .X(_3360_));
 sky130_fd_sc_hd__clkbuf_1 _8214_ (.A(_3360_),
    .X(_0040_));
 sky130_fd_sc_hd__and2_1 _8215_ (.A(_3357_),
    .B(net63),
    .X(_3361_));
 sky130_fd_sc_hd__clkbuf_1 _8216_ (.A(_3361_),
    .X(_0041_));
 sky130_fd_sc_hd__and2_1 _8217_ (.A(_3357_),
    .B(net64),
    .X(_3363_));
 sky130_fd_sc_hd__clkbuf_1 _8218_ (.A(_3363_),
    .X(_0042_));
 sky130_fd_sc_hd__and2_1 _8219_ (.A(_3357_),
    .B(net34),
    .X(_3364_));
 sky130_fd_sc_hd__clkbuf_1 _8220_ (.A(_3364_),
    .X(_0043_));
 sky130_fd_sc_hd__and2_1 _8221_ (.A(_3357_),
    .B(net35),
    .X(_3365_));
 sky130_fd_sc_hd__clkbuf_1 _8222_ (.A(_3365_),
    .X(_0044_));
 sky130_fd_sc_hd__and2_1 _8223_ (.A(_3357_),
    .B(net36),
    .X(_3366_));
 sky130_fd_sc_hd__clkbuf_1 _8224_ (.A(_3366_),
    .X(_0045_));
 sky130_fd_sc_hd__and2_1 _8225_ (.A(_3357_),
    .B(net37),
    .X(_3367_));
 sky130_fd_sc_hd__clkbuf_1 _8226_ (.A(_3367_),
    .X(_0046_));
 sky130_fd_sc_hd__and2_1 _8227_ (.A(_3357_),
    .B(net38),
    .X(_3369_));
 sky130_fd_sc_hd__clkbuf_1 _8228_ (.A(_3369_),
    .X(_0047_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _8229_ (.A(net65),
    .X(_3370_));
 sky130_fd_sc_hd__and2_1 _8230_ (.A(_3370_),
    .B(net39),
    .X(_3371_));
 sky130_fd_sc_hd__clkbuf_1 _8231_ (.A(_3371_),
    .X(_0048_));
 sky130_fd_sc_hd__and2_1 _8232_ (.A(_3370_),
    .B(net40),
    .X(_3372_));
 sky130_fd_sc_hd__clkbuf_1 _8233_ (.A(_3372_),
    .X(_0049_));
 sky130_fd_sc_hd__and2_1 _8234_ (.A(_3370_),
    .B(net41),
    .X(_3373_));
 sky130_fd_sc_hd__clkbuf_1 _8235_ (.A(_3373_),
    .X(_0050_));
 sky130_fd_sc_hd__and2_1 _8236_ (.A(_3370_),
    .B(net42),
    .X(_3375_));
 sky130_fd_sc_hd__clkbuf_1 _8237_ (.A(_3375_),
    .X(_0051_));
 sky130_fd_sc_hd__and2_1 _8238_ (.A(_3370_),
    .B(net43),
    .X(_3376_));
 sky130_fd_sc_hd__clkbuf_1 _8239_ (.A(_3376_),
    .X(_0052_));
 sky130_fd_sc_hd__and2_1 _8240_ (.A(_3370_),
    .B(net45),
    .X(_3377_));
 sky130_fd_sc_hd__clkbuf_1 _8241_ (.A(_3377_),
    .X(_0053_));
 sky130_fd_sc_hd__and2_1 _8242_ (.A(_3370_),
    .B(net46),
    .X(_3378_));
 sky130_fd_sc_hd__clkbuf_1 _8243_ (.A(_3378_),
    .X(_0054_));
 sky130_fd_sc_hd__and2_1 _8244_ (.A(_3370_),
    .B(net47),
    .X(_3379_));
 sky130_fd_sc_hd__buf_1 _8245_ (.A(_3379_),
    .X(_0055_));
 sky130_fd_sc_hd__and2_1 _8246_ (.A(_3370_),
    .B(net48),
    .X(_3381_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _8247_ (.A(_3381_),
    .X(_0056_));
 sky130_fd_sc_hd__and2_1 _8248_ (.A(_3370_),
    .B(net49),
    .X(_3382_));
 sky130_fd_sc_hd__buf_1 _8249_ (.A(_3382_),
    .X(_0057_));
 sky130_fd_sc_hd__buf_2 _8250_ (.A(net65),
    .X(_3383_));
 sky130_fd_sc_hd__and2_1 _8251_ (.A(_3383_),
    .B(net50),
    .X(_3384_));
 sky130_fd_sc_hd__clkbuf_1 _8252_ (.A(_3384_),
    .X(_0058_));
 sky130_fd_sc_hd__and2_1 _8253_ (.A(_3383_),
    .B(net51),
    .X(_3385_));
 sky130_fd_sc_hd__clkbuf_1 _8254_ (.A(_3385_),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _8255_ (.A(_3383_),
    .B(net52),
    .X(_3386_));
 sky130_fd_sc_hd__clkbuf_1 _8256_ (.A(_3386_),
    .X(_0060_));
 sky130_fd_sc_hd__and2_1 _8257_ (.A(_3383_),
    .B(net53),
    .X(_3388_));
 sky130_fd_sc_hd__clkbuf_1 _8258_ (.A(_3388_),
    .X(_0061_));
 sky130_fd_sc_hd__and2_1 _8259_ (.A(_3383_),
    .B(net54),
    .X(_3389_));
 sky130_fd_sc_hd__clkbuf_1 _8260_ (.A(_3389_),
    .X(_0062_));
 sky130_fd_sc_hd__and2_1 _8261_ (.A(_3383_),
    .B(net56),
    .X(_3390_));
 sky130_fd_sc_hd__clkbuf_1 _8262_ (.A(_3390_),
    .X(_0063_));
 sky130_fd_sc_hd__and2_1 _8263_ (.A(_3383_),
    .B(net57),
    .X(_3391_));
 sky130_fd_sc_hd__clkbuf_1 _8264_ (.A(_3391_),
    .X(_0064_));
 sky130_fd_sc_hd__inv_2 _8265_ (.A(_2752_),
    .Y(_3392_));
 sky130_fd_sc_hd__inv_2 _8266_ (.A(_2767_),
    .Y(_3394_));
 sky130_fd_sc_hd__nor2_1 _8267_ (.A(_3394_),
    .B(_2790_),
    .Y(_3395_));
 sky130_fd_sc_hd__inv_2 _8268_ (.A(_2801_),
    .Y(_3396_));
 sky130_fd_sc_hd__nor2_1 _8269_ (.A(_3396_),
    .B(_2813_),
    .Y(_3397_));
 sky130_fd_sc_hd__a21o_1 _8270_ (.A1(_2816_),
    .A2(_3395_),
    .B1(_3397_),
    .X(_3398_));
 sky130_fd_sc_hd__inv_2 _8271_ (.A(_2723_),
    .Y(_3399_));
 sky130_fd_sc_hd__nor2_1 _8272_ (.A(_3399_),
    .B(_2749_),
    .Y(_3400_));
 sky130_fd_sc_hd__xnor2_2 _8273_ (.A(\F1.sign_b ),
    .B(_3346_),
    .Y(_3401_));
 sky130_fd_sc_hd__a211o_1 _8274_ (.A1(_3392_),
    .A2(_3398_),
    .B1(_3400_),
    .C1(_3401_),
    .X(_3402_));
 sky130_fd_sc_hd__or2_1 _8275_ (.A(net119),
    .B(_3402_),
    .X(_3403_));
 sky130_fd_sc_hd__inv_2 _8276_ (.A(_3403_),
    .Y(_3405_));
 sky130_fd_sc_hd__inv_2 _8277_ (.A(_3276_),
    .Y(_3406_));
 sky130_fd_sc_hd__nor2_1 _8278_ (.A(_3406_),
    .B(_3279_),
    .Y(_3407_));
 sky130_fd_sc_hd__nand2_2 _8279_ (.A(_3273_),
    .B(_3280_),
    .Y(_3408_));
 sky130_fd_sc_hd__or3_4 _8280_ (.A(_3287_),
    .B(_3293_),
    .C(_3408_),
    .X(_3409_));
 sky130_fd_sc_hd__inv_2 _8281_ (.A(_3248_),
    .Y(_3410_));
 sky130_fd_sc_hd__nor2_1 _8282_ (.A(_3410_),
    .B(_3252_),
    .Y(_3411_));
 sky130_fd_sc_hd__inv_2 _8283_ (.A(_3258_),
    .Y(_3412_));
 sky130_fd_sc_hd__nor2_1 _8284_ (.A(_3412_),
    .B(_3262_),
    .Y(_3413_));
 sky130_fd_sc_hd__a21o_1 _8285_ (.A1(_3265_),
    .A2(_3411_),
    .B1(_3413_),
    .X(_3414_));
 sky130_fd_sc_hd__and2_1 _8286_ (.A(_3303_),
    .B(_3311_),
    .X(_3416_));
 sky130_fd_sc_hd__inv_2 _8287_ (.A(_3307_),
    .Y(_3417_));
 sky130_fd_sc_hd__nor2_1 _8288_ (.A(_3417_),
    .B(_3310_),
    .Y(_3418_));
 sky130_fd_sc_hd__inv_2 _8289_ (.A(_3299_),
    .Y(_3419_));
 sky130_fd_sc_hd__nor2_1 _8290_ (.A(_3419_),
    .B(_3302_),
    .Y(_3420_));
 sky130_fd_sc_hd__a21o_1 _8291_ (.A1(net116),
    .A2(_3418_),
    .B1(_3420_),
    .X(_3421_));
 sky130_fd_sc_hd__a21oi_1 _8292_ (.A1(_3414_),
    .A2(_3416_),
    .B1(_3421_),
    .Y(_3422_));
 sky130_fd_sc_hd__inv_2 _8293_ (.A(_3284_),
    .Y(_3423_));
 sky130_fd_sc_hd__or2_1 _8294_ (.A(_3423_),
    .B(_3286_),
    .X(_3424_));
 sky130_fd_sc_hd__inv_2 _8295_ (.A(_3292_),
    .Y(_3425_));
 sky130_fd_sc_hd__nand2_1 _8296_ (.A(_3289_),
    .B(_3425_),
    .Y(_3427_));
 sky130_fd_sc_hd__o21a_1 _8297_ (.A1(_3293_),
    .A2(_3424_),
    .B1(_3427_),
    .X(_3428_));
 sky130_fd_sc_hd__nand2_1 _8298_ (.A(_3269_),
    .B(_3271_),
    .Y(_3429_));
 sky130_fd_sc_hd__o221a_1 _8299_ (.A1(_3409_),
    .A2(_3422_),
    .B1(_3428_),
    .B2(_3408_),
    .C1(_3429_),
    .X(_3430_));
 sky130_fd_sc_hd__a21boi_1 _8300_ (.A1(_3273_),
    .A2(_3407_),
    .B1_N(_3430_),
    .Y(_3431_));
 sky130_fd_sc_hd__inv_2 _8301_ (.A(_2954_),
    .Y(_3432_));
 sky130_fd_sc_hd__nor2_1 _8302_ (.A(_3432_),
    .B(_3009_),
    .Y(_3433_));
 sky130_fd_sc_hd__nand2_1 _8303_ (.A(_3094_),
    .B(_3095_),
    .Y(_3434_));
 sky130_fd_sc_hd__nand2_1 _8304_ (.A(_3125_),
    .B(_3126_),
    .Y(_3435_));
 sky130_fd_sc_hd__or2_4 _8305_ (.A(_3010_),
    .B(_3060_),
    .X(_3436_));
 sky130_fd_sc_hd__inv_2 _8306_ (.A(_3436_),
    .Y(_3438_));
 sky130_fd_sc_hd__or2_1 _8307_ (.A(_3139_),
    .B(_3153_),
    .X(_3439_));
 sky130_fd_sc_hd__nand2_1 _8308_ (.A(_3235_),
    .B(_3439_),
    .Y(_3440_));
 sky130_fd_sc_hd__and3_1 _8309_ (.A(_3212_),
    .B(_3220_),
    .C(_3231_),
    .X(_3441_));
 sky130_fd_sc_hd__nor2_2 _8310_ (.A(_3233_),
    .B(_3441_),
    .Y(_3442_));
 sky130_fd_sc_hd__xnor2_2 _8311_ (.A(_3182_),
    .B(net112),
    .Y(_3443_));
 sky130_fd_sc_hd__o21ba_1 _8312_ (.A1(_3185_),
    .A2(_3196_),
    .B1_N(_3210_),
    .X(_3444_));
 sky130_fd_sc_hd__a21o_1 _8313_ (.A1(_2844_),
    .A2(_3179_),
    .B1(_3181_),
    .X(_3445_));
 sky130_fd_sc_hd__nand2_1 _8314_ (.A(_3165_),
    .B(_3445_),
    .Y(_3446_));
 sky130_fd_sc_hd__a21boi_1 _8315_ (.A1(_3443_),
    .A2(_3444_),
    .B1_N(_3446_),
    .Y(_3447_));
 sky130_fd_sc_hd__a21bo_1 _8316_ (.A1(_3212_),
    .A2(_3220_),
    .B1_N(_3231_),
    .X(_3449_));
 sky130_fd_sc_hd__o21ai_1 _8317_ (.A1(_3447_),
    .A2(_3442_),
    .B1(_3449_),
    .Y(_3450_));
 sky130_fd_sc_hd__inv_2 _8318_ (.A(_3139_),
    .Y(_3451_));
 sky130_fd_sc_hd__nor2_1 _8319_ (.A(_3451_),
    .B(_3153_),
    .Y(_3452_));
 sky130_fd_sc_hd__a21o_1 _8320_ (.A1(_3450_),
    .A2(_3440_),
    .B1(_3452_),
    .X(_3453_));
 sky130_fd_sc_hd__o2bb2a_1 _8321_ (.A1_N(_3061_),
    .A2_N(_3076_),
    .B1(_3080_),
    .B2(_3093_),
    .X(_3454_));
 sky130_fd_sc_hd__a21boi_1 _8322_ (.A1(_3110_),
    .A2(_3124_),
    .B1_N(_3109_),
    .Y(_3455_));
 sky130_fd_sc_hd__a21oi_1 _8323_ (.A1(_3435_),
    .A2(_3454_),
    .B1(_3455_),
    .Y(_3456_));
 sky130_fd_sc_hd__nor2_1 _8324_ (.A(_3029_),
    .B(_3059_),
    .Y(_3457_));
 sky130_fd_sc_hd__and2b_1 _8325_ (.A_N(_3010_),
    .B(_3457_),
    .X(_3458_));
 sky130_fd_sc_hd__o21bai_1 _8326_ (.A1(_3436_),
    .A2(_3456_),
    .B1_N(_3458_),
    .Y(_3460_));
 sky130_fd_sc_hd__a41o_1 _8327_ (.A1(_3453_),
    .A2(_3435_),
    .A3(_3438_),
    .A4(_3434_),
    .B1(_3460_),
    .X(_3461_));
 sky130_fd_sc_hd__and3b_1 _8328_ (.A_N(_3409_),
    .B(_3265_),
    .C(_3255_),
    .X(_3462_));
 sky130_fd_sc_hd__o211ai_2 _8329_ (.A1(_3433_),
    .A2(_3461_),
    .B1(_3462_),
    .C1(_3416_),
    .Y(_3463_));
 sky130_fd_sc_hd__inv_2 _8330_ (.A(_2904_),
    .Y(_3464_));
 sky130_fd_sc_hd__inv_2 _8331_ (.A(_2932_),
    .Y(_3465_));
 sky130_fd_sc_hd__nand2_1 _8332_ (.A(_2848_),
    .B(_2877_),
    .Y(_3466_));
 sky130_fd_sc_hd__a2111o_1 _8333_ (.A1(_3463_),
    .A2(_3431_),
    .B1(_3464_),
    .C1(_3465_),
    .D1(_3466_),
    .X(_3467_));
 sky130_fd_sc_hd__nand2_1 _8334_ (.A(_2928_),
    .B(_2922_),
    .Y(_3468_));
 sky130_fd_sc_hd__nand2_1 _8335_ (.A(_2901_),
    .B(_2893_),
    .Y(_3469_));
 sky130_fd_sc_hd__o21a_1 _8336_ (.A1(_3464_),
    .A2(_3468_),
    .B1(_3469_),
    .X(_3471_));
 sky130_fd_sc_hd__inv_2 _8337_ (.A(_2859_),
    .Y(_3472_));
 sky130_fd_sc_hd__nor2_1 _8338_ (.A(_3472_),
    .B(_2873_),
    .Y(_3473_));
 sky130_fd_sc_hd__and2b_1 _8339_ (.A_N(_2829_),
    .B(_2845_),
    .X(_3474_));
 sky130_fd_sc_hd__a21oi_1 _8340_ (.A1(_2848_),
    .A2(_3473_),
    .B1(_3474_),
    .Y(_3475_));
 sky130_fd_sc_hd__o21a_1 _8341_ (.A1(_3466_),
    .A2(_3471_),
    .B1(_3475_),
    .X(_3476_));
 sky130_fd_sc_hd__and2_1 _8342_ (.A(_3392_),
    .B(_2816_),
    .X(_3477_));
 sky130_fd_sc_hd__inv_2 _8343_ (.A(_3477_),
    .Y(_3478_));
 sky130_fd_sc_hd__inv_2 _8344_ (.A(_2793_),
    .Y(_3479_));
 sky130_fd_sc_hd__a211o_4 _8345_ (.A1(_3476_),
    .A2(_3467_),
    .B1(_3478_),
    .C1(_3479_),
    .X(_3480_));
 sky130_fd_sc_hd__a21oi_4 _8346_ (.A1(_3480_),
    .A2(_3405_),
    .B1(_3401_),
    .Y(_3482_));
 sky130_fd_sc_hd__or2b_4 _8347_ (.A(_3402_),
    .B_N(_3480_),
    .X(_3483_));
 sky130_fd_sc_hd__o21ai_4 _8348_ (.A1(_2818_),
    .A2(net102),
    .B1(_3343_),
    .Y(_3484_));
 sky130_fd_sc_hd__xor2_1 _8349_ (.A(\F1.sign_b ),
    .B(_3346_),
    .X(_3485_));
 sky130_fd_sc_hd__clkbuf_4 _8350_ (.A(_3485_),
    .X(_3486_));
 sky130_fd_sc_hd__inv_2 _8351_ (.A(_2792_),
    .Y(_3487_));
 sky130_fd_sc_hd__a21oi_1 _8352_ (.A1(_2815_),
    .A2(_3487_),
    .B1(_2814_),
    .Y(_3488_));
 sky130_fd_sc_hd__o211a_1 _8353_ (.A1(_2818_),
    .A2(net104),
    .B1(_3488_),
    .C1(_3343_),
    .X(_3489_));
 sky130_fd_sc_hd__a211o_1 _8354_ (.A1(_3340_),
    .A2(_3484_),
    .B1(_3486_),
    .C1(_3489_),
    .X(_3490_));
 sky130_fd_sc_hd__o21a_1 _8355_ (.A1(_3185_),
    .A2(_3196_),
    .B1(_3210_),
    .X(_3491_));
 sky130_fd_sc_hd__and2_1 _8356_ (.A(_3165_),
    .B(_3182_),
    .X(_3493_));
 sky130_fd_sc_hd__a211oi_2 _8357_ (.A1(_3183_),
    .A2(_3491_),
    .B1(_3233_),
    .C1(_3493_),
    .Y(_3494_));
 sky130_fd_sc_hd__o31ai_2 _8358_ (.A1(_3154_),
    .A2(_3441_),
    .A3(_3494_),
    .B1(_3235_),
    .Y(_3495_));
 sky130_fd_sc_hd__nand2_1 _8359_ (.A(_3126_),
    .B(_3095_),
    .Y(_3496_));
 sky130_fd_sc_hd__nand4_1 _8360_ (.A(_3010_),
    .B(_3060_),
    .C(_3125_),
    .D(_3496_),
    .Y(_3497_));
 sky130_fd_sc_hd__or2_1 _8361_ (.A(_3242_),
    .B(_3059_),
    .X(_3498_));
 sky130_fd_sc_hd__a21o_1 _8362_ (.A1(_3240_),
    .A2(_3498_),
    .B1(_3237_),
    .X(_3499_));
 sky130_fd_sc_hd__o211ai_2 _8363_ (.A1(_3128_),
    .A2(_3495_),
    .B1(_3497_),
    .C1(_3499_),
    .Y(_3500_));
 sky130_fd_sc_hd__a21boi_1 _8364_ (.A1(_3254_),
    .A2(_3264_),
    .B1_N(_3263_),
    .Y(_3501_));
 sky130_fd_sc_hd__nor2_1 _8365_ (.A(_3307_),
    .B(_3310_),
    .Y(_3502_));
 sky130_fd_sc_hd__o21ai_1 _8366_ (.A1(_3317_),
    .A2(_3502_),
    .B1(_3314_),
    .Y(_3504_));
 sky130_fd_sc_hd__a21bo_1 _8367_ (.A1(_3312_),
    .A2(_3501_),
    .B1_N(_3504_),
    .X(_3505_));
 sky130_fd_sc_hd__or2_1 _8368_ (.A(_3276_),
    .B(_3279_),
    .X(_3506_));
 sky130_fd_sc_hd__o21ai_1 _8369_ (.A1(_3326_),
    .A2(_3506_),
    .B1(_3324_),
    .Y(_3507_));
 sky130_fd_sc_hd__nor2_1 _8370_ (.A(_3284_),
    .B(_3286_),
    .Y(_3508_));
 sky130_fd_sc_hd__o211a_1 _8371_ (.A1(_3508_),
    .A2(_3322_),
    .B1(_3321_),
    .C1(_3319_),
    .X(_3509_));
 sky130_fd_sc_hd__a211o_1 _8372_ (.A1(_3296_),
    .A2(_3505_),
    .B1(_3507_),
    .C1(_3509_),
    .X(_3510_));
 sky130_fd_sc_hd__a21o_1 _8373_ (.A1(_3313_),
    .A2(_3500_),
    .B1(_3510_),
    .X(_3511_));
 sky130_fd_sc_hd__nand2_1 _8374_ (.A(_2847_),
    .B(_2875_),
    .Y(_3512_));
 sky130_fd_sc_hd__a21o_1 _8375_ (.A1(_2903_),
    .A2(_2930_),
    .B1(_2902_),
    .X(_3513_));
 sky130_fd_sc_hd__inv_2 _8376_ (.A(_3513_),
    .Y(_3515_));
 sky130_fd_sc_hd__a22o_1 _8377_ (.A1(_2846_),
    .A2(_3512_),
    .B1(_2878_),
    .B2(_3515_),
    .X(_3516_));
 sky130_fd_sc_hd__a21oi_1 _8378_ (.A1(_2934_),
    .A2(_3511_),
    .B1(_3516_),
    .Y(_3517_));
 sky130_fd_sc_hd__o211a_1 _8379_ (.A1(_2818_),
    .A2(net102),
    .B1(_3517_),
    .C1(_3343_),
    .X(_3518_));
 sky130_fd_sc_hd__a2111o_1 _8380_ (.A1(_3484_),
    .A2(net103),
    .B1(_3485_),
    .C1(_3518_),
    .D1(_2817_),
    .X(_3519_));
 sky130_fd_sc_hd__a21o_1 _8381_ (.A1(_3519_),
    .A2(_3490_),
    .B1(_3392_),
    .X(_3520_));
 sky130_fd_sc_hd__a21o_1 _8382_ (.A1(_2661_),
    .A2(_2751_),
    .B1(_3341_),
    .X(_3521_));
 sky130_fd_sc_hd__and2_1 _8383_ (.A(_3401_),
    .B(_3521_),
    .X(_3522_));
 sky130_fd_sc_hd__inv_2 _8384_ (.A(_3522_),
    .Y(_3523_));
 sky130_fd_sc_hd__a31o_4 _8385_ (.A1(_3520_),
    .A2(_3483_),
    .A3(_3523_),
    .B1(net119),
    .X(_3524_));
 sky130_fd_sc_hd__nand4_2 _8386_ (.A(_3520_),
    .B(_3483_),
    .C(net120),
    .D(_3523_),
    .Y(_3526_));
 sky130_fd_sc_hd__nand2_4 _8387_ (.A(_3524_),
    .B(_3526_),
    .Y(_3527_));
 sky130_fd_sc_hd__or2_4 _8388_ (.A(_3482_),
    .B(_3527_),
    .X(_3528_));
 sky130_fd_sc_hd__buf_6 _8389_ (.A(_3528_),
    .X(_3529_));
 sky130_fd_sc_hd__buf_4 _8390_ (.A(_3529_),
    .X(_3530_));
 sky130_fd_sc_hd__or3_1 _8391_ (.A(_3185_),
    .B(_3196_),
    .C(_3210_),
    .X(_3531_));
 sky130_fd_sc_hd__inv_2 _8392_ (.A(_3491_),
    .Y(_3532_));
 sky130_fd_sc_hd__nand2_1 _8393_ (.A(_3531_),
    .B(_3532_),
    .Y(_3533_));
 sky130_fd_sc_hd__clkbuf_4 _8394_ (.A(_3401_),
    .X(_3534_));
 sky130_fd_sc_hd__clkbuf_4 _8395_ (.A(_3534_),
    .X(_3535_));
 sky130_fd_sc_hd__mux2_1 _8396_ (.A0(_3531_),
    .A1(_3532_),
    .S(_3345_),
    .X(_3537_));
 sky130_fd_sc_hd__nor2_1 _8397_ (.A(_3535_),
    .B(_3444_),
    .Y(_3538_));
 sky130_fd_sc_hd__a21oi_1 _8398_ (.A1(_3535_),
    .A2(_3537_),
    .B1(_3538_),
    .Y(_3539_));
 sky130_fd_sc_hd__xor2_1 _8399_ (.A(_3443_),
    .B(_3539_),
    .X(_3540_));
 sky130_fd_sc_hd__mux2_1 _8400_ (.A0(_3533_),
    .A1(_3540_),
    .S(net111),
    .X(_3541_));
 sky130_fd_sc_hd__and3_1 _8401_ (.A(_3348_),
    .B(_3530_),
    .C(_3541_),
    .X(_3542_));
 sky130_fd_sc_hd__clkbuf_1 _8402_ (.A(_3542_),
    .X(_0065_));
 sky130_fd_sc_hd__buf_2 _8403_ (.A(_3524_),
    .X(_3543_));
 sky130_fd_sc_hd__buf_2 _8404_ (.A(net111),
    .X(_3544_));
 sky130_fd_sc_hd__and2_1 _8405_ (.A(_3183_),
    .B(_3211_),
    .X(_3545_));
 sky130_fd_sc_hd__a21oi_1 _8406_ (.A1(_3183_),
    .A2(_3491_),
    .B1(_3493_),
    .Y(_3547_));
 sky130_fd_sc_hd__mux2_1 _8407_ (.A0(_3545_),
    .A1(_3547_),
    .S(_3345_),
    .X(_3548_));
 sky130_fd_sc_hd__mux2_1 _8408_ (.A0(_3447_),
    .A1(_3548_),
    .S(_3535_),
    .X(_3549_));
 sky130_fd_sc_hd__xnor2_1 _8409_ (.A(_3442_),
    .B(_3549_),
    .Y(_3550_));
 sky130_fd_sc_hd__nand2_1 _8410_ (.A(_3544_),
    .B(_3550_),
    .Y(_3551_));
 sky130_fd_sc_hd__o211a_1 _8411_ (.A1(net133),
    .A2(_3533_),
    .B1(_3551_),
    .C1(_3383_),
    .X(_3552_));
 sky130_fd_sc_hd__o21a_1 _8412_ (.A1(_3543_),
    .A2(_3540_),
    .B1(_3552_),
    .X(_0066_));
 sky130_fd_sc_hd__a31oi_4 _8413_ (.A1(_3483_),
    .A2(_3520_),
    .A3(_3523_),
    .B1(net121),
    .Y(_3553_));
 sky130_fd_sc_hd__nor2_1 _8414_ (.A(_3441_),
    .B(_3494_),
    .Y(_3554_));
 sky130_fd_sc_hd__mux2_1 _8415_ (.A0(_3234_),
    .A1(_3554_),
    .S(_3345_),
    .X(_3555_));
 sky130_fd_sc_hd__mux2_1 _8416_ (.A0(_3450_),
    .A1(_3555_),
    .S(_3535_),
    .X(_3557_));
 sky130_fd_sc_hd__xor2_1 _8417_ (.A(_3440_),
    .B(_3557_),
    .X(_3558_));
 sky130_fd_sc_hd__a21o_1 _8418_ (.A1(_3405_),
    .A2(_3480_),
    .B1(_3534_),
    .X(_3559_));
 sky130_fd_sc_hd__buf_2 _8419_ (.A(_3559_),
    .X(_3560_));
 sky130_fd_sc_hd__o2bb2a_1 _8420_ (.A1_N(_3553_),
    .A2_N(_3550_),
    .B1(_3558_),
    .B2(_3560_),
    .X(_3561_));
 sky130_fd_sc_hd__o211a_1 _8421_ (.A1(_3530_),
    .A2(_3540_),
    .B1(_3561_),
    .C1(_3350_),
    .X(_0067_));
 sky130_fd_sc_hd__and3_1 _8422_ (.A(_3559_),
    .B(_3524_),
    .C(_3526_),
    .X(_3562_));
 sky130_fd_sc_hd__buf_2 _8423_ (.A(_3562_),
    .X(_3563_));
 sky130_fd_sc_hd__mux2_2 _8424_ (.A0(_3236_),
    .A1(_3495_),
    .S(_3344_),
    .X(_3564_));
 sky130_fd_sc_hd__mux2_1 _8425_ (.A0(_3453_),
    .A1(_3564_),
    .S(_3535_),
    .X(_3565_));
 sky130_fd_sc_hd__xnor2_1 _8426_ (.A(_3097_),
    .B(_3565_),
    .Y(_3567_));
 sky130_fd_sc_hd__o221a_1 _8427_ (.A1(_3543_),
    .A2(_3558_),
    .B1(_3567_),
    .B2(_3560_),
    .C1(_3348_),
    .X(_3568_));
 sky130_fd_sc_hd__a21boi_1 _8428_ (.A1(_3563_),
    .A2(_3550_),
    .B1_N(_3568_),
    .Y(_0068_));
 sky130_fd_sc_hd__clkbuf_4 _8429_ (.A(_3534_),
    .X(_3569_));
 sky130_fd_sc_hd__or2_1 _8430_ (.A(_3434_),
    .B(_3564_),
    .X(_3570_));
 sky130_fd_sc_hd__mux2_1 _8431_ (.A0(_3094_),
    .A1(_3095_),
    .S(_3345_),
    .X(_3571_));
 sky130_fd_sc_hd__and2_1 _8432_ (.A(_3434_),
    .B(_3453_),
    .X(_3572_));
 sky130_fd_sc_hd__o21a_1 _8433_ (.A1(_3572_),
    .A2(_3454_),
    .B1(_3486_),
    .X(_3573_));
 sky130_fd_sc_hd__a31o_1 _8434_ (.A1(_3569_),
    .A2(_3570_),
    .A3(_3571_),
    .B1(_3573_),
    .X(_3574_));
 sky130_fd_sc_hd__xnor2_1 _8435_ (.A(_3127_),
    .B(_3574_),
    .Y(_3575_));
 sky130_fd_sc_hd__o221a_1 _8436_ (.A1(_3543_),
    .A2(_3567_),
    .B1(_3575_),
    .B2(_3560_),
    .C1(_3348_),
    .X(_3577_));
 sky130_fd_sc_hd__o21a_1 _8437_ (.A1(_3530_),
    .A2(_3558_),
    .B1(_3577_),
    .X(_0069_));
 sky130_fd_sc_hd__inv_2 _8438_ (.A(_3060_),
    .Y(_3578_));
 sky130_fd_sc_hd__a21bo_1 _8439_ (.A1(_3435_),
    .A2(_3572_),
    .B1_N(_3456_),
    .X(_3579_));
 sky130_fd_sc_hd__nand2_1 _8440_ (.A(_3125_),
    .B(_3496_),
    .Y(_3580_));
 sky130_fd_sc_hd__mux2_1 _8441_ (.A0(_3238_),
    .A1(_3580_),
    .S(_3344_),
    .X(_3581_));
 sky130_fd_sc_hd__o31a_1 _8442_ (.A1(_3434_),
    .A2(_3435_),
    .A3(_3564_),
    .B1(_3581_),
    .X(_3582_));
 sky130_fd_sc_hd__mux2_1 _8443_ (.A0(_3579_),
    .A1(_3582_),
    .S(_3535_),
    .X(_3583_));
 sky130_fd_sc_hd__xnor2_2 _8444_ (.A(_3578_),
    .B(_3583_),
    .Y(_3584_));
 sky130_fd_sc_hd__nor2_1 _8445_ (.A(_3559_),
    .B(_3584_),
    .Y(_3585_));
 sky130_fd_sc_hd__a211o_1 _8446_ (.A1(_3560_),
    .A2(_3575_),
    .B1(_3585_),
    .C1(_3563_),
    .X(_3587_));
 sky130_fd_sc_hd__o211a_1 _8447_ (.A1(_3530_),
    .A2(_3567_),
    .B1(_3587_),
    .C1(_3350_),
    .X(_0070_));
 sky130_fd_sc_hd__a21o_1 _8448_ (.A1(_3578_),
    .A2(_3579_),
    .B1(_3457_),
    .X(_3588_));
 sky130_fd_sc_hd__buf_4 _8449_ (.A(_3484_),
    .X(_3589_));
 sky130_fd_sc_hd__nand2_1 _8450_ (.A(_3243_),
    .B(_3589_),
    .Y(_3590_));
 sky130_fd_sc_hd__o21a_1 _8451_ (.A1(_3498_),
    .A2(_3589_),
    .B1(_3590_),
    .X(_3591_));
 sky130_fd_sc_hd__o211a_1 _8452_ (.A1(_3578_),
    .A2(_3582_),
    .B1(_3591_),
    .C1(_3535_),
    .X(_3592_));
 sky130_fd_sc_hd__a21oi_1 _8453_ (.A1(_3486_),
    .A2(_3588_),
    .B1(_3592_),
    .Y(_3593_));
 sky130_fd_sc_hd__xnor2_1 _8454_ (.A(_3010_),
    .B(_3593_),
    .Y(_3594_));
 sky130_fd_sc_hd__a2bb2o_1 _8455_ (.A1_N(_3529_),
    .A2_N(_3575_),
    .B1(_3584_),
    .B2(_3553_),
    .X(_3595_));
 sky130_fd_sc_hd__inv_2 _8456_ (.A(net65),
    .Y(_3597_));
 sky130_fd_sc_hd__a211oi_1 _8457_ (.A1(_3544_),
    .A2(_3594_),
    .B1(_3595_),
    .C1(_3597_),
    .Y(_0071_));
 sky130_fd_sc_hd__nor2_1 _8458_ (.A(_3433_),
    .B(_3461_),
    .Y(_3598_));
 sky130_fd_sc_hd__mux2_4 _8459_ (.A0(_3245_),
    .A1(_3500_),
    .S(_3344_),
    .X(_3599_));
 sky130_fd_sc_hd__mux2_1 _8460_ (.A0(_3598_),
    .A1(_3599_),
    .S(_3534_),
    .X(_3600_));
 sky130_fd_sc_hd__xnor2_2 _8461_ (.A(_3255_),
    .B(_3600_),
    .Y(_3601_));
 sky130_fd_sc_hd__inv_2 _8462_ (.A(_3601_),
    .Y(_3602_));
 sky130_fd_sc_hd__a221o_1 _8463_ (.A1(_3553_),
    .A2(_3594_),
    .B1(_3602_),
    .B2(_3544_),
    .C1(_3597_),
    .X(_3603_));
 sky130_fd_sc_hd__a21oi_1 _8464_ (.A1(_3563_),
    .A2(_3584_),
    .B1(_3603_),
    .Y(_0072_));
 sky130_fd_sc_hd__nor2_1 _8465_ (.A(_3253_),
    .B(_3344_),
    .Y(_3604_));
 sky130_fd_sc_hd__nor2_1 _8466_ (.A(_3254_),
    .B(_3484_),
    .Y(_3606_));
 sky130_fd_sc_hd__a311o_1 _8467_ (.A1(_3253_),
    .A2(_3254_),
    .A3(_3599_),
    .B1(_3604_),
    .C1(_3606_),
    .X(_3607_));
 sky130_fd_sc_hd__or3_1 _8468_ (.A(_3438_),
    .B(_3458_),
    .C(_3433_),
    .X(_3608_));
 sky130_fd_sc_hd__or3b_1 _8469_ (.A(_3458_),
    .B(_3433_),
    .C_N(_3456_),
    .X(_3609_));
 sky130_fd_sc_hd__a31o_1 _8470_ (.A1(_3434_),
    .A2(_3435_),
    .A3(_3453_),
    .B1(_3609_),
    .X(_3610_));
 sky130_fd_sc_hd__a31oi_1 _8471_ (.A1(_3255_),
    .A2(_3608_),
    .A3(_3610_),
    .B1(_3411_),
    .Y(_3611_));
 sky130_fd_sc_hd__mux2_2 _8472_ (.A0(_3607_),
    .A1(_3611_),
    .S(_3486_),
    .X(_3612_));
 sky130_fd_sc_hd__xor2_2 _8473_ (.A(_3265_),
    .B(_3612_),
    .X(_3613_));
 sky130_fd_sc_hd__mux2_4 _8474_ (.A0(_3602_),
    .A1(_3613_),
    .S(_3482_),
    .X(_3614_));
 sky130_fd_sc_hd__mux2_1 _8475_ (.A0(_3594_),
    .A1(_3614_),
    .S(_3529_),
    .X(_3615_));
 sky130_fd_sc_hd__nor2_1 _8476_ (.A(_3597_),
    .B(_3615_),
    .Y(_0073_));
 sky130_fd_sc_hd__nand2_1 _8477_ (.A(_3559_),
    .B(_3613_),
    .Y(_3617_));
 sky130_fd_sc_hd__nand2_1 _8478_ (.A(_3245_),
    .B(_3266_),
    .Y(_3618_));
 sky130_fd_sc_hd__a21oi_1 _8479_ (.A1(_3266_),
    .A2(_3500_),
    .B1(_3501_),
    .Y(_3619_));
 sky130_fd_sc_hd__o211a_1 _8480_ (.A1(_2818_),
    .A2(_3339_),
    .B1(_3619_),
    .C1(_3343_),
    .X(_3620_));
 sky130_fd_sc_hd__a31o_1 _8481_ (.A1(_3330_),
    .A2(_3484_),
    .A3(_3618_),
    .B1(_3620_),
    .X(_3621_));
 sky130_fd_sc_hd__a41o_1 _8482_ (.A1(_3255_),
    .A2(_3265_),
    .A3(_3608_),
    .A4(_3610_),
    .B1(_3414_),
    .X(_3622_));
 sky130_fd_sc_hd__and2_1 _8483_ (.A(_3486_),
    .B(_3622_),
    .X(_3623_));
 sky130_fd_sc_hd__a21o_1 _8484_ (.A1(_3569_),
    .A2(_3621_),
    .B1(_3623_),
    .X(_3624_));
 sky130_fd_sc_hd__xnor2_2 _8485_ (.A(_3311_),
    .B(_3624_),
    .Y(_3625_));
 sky130_fd_sc_hd__nand2_1 _8486_ (.A(_3544_),
    .B(_3625_),
    .Y(_3627_));
 sky130_fd_sc_hd__a21o_1 _8487_ (.A1(_3617_),
    .A2(_3627_),
    .B1(_3563_),
    .X(_3628_));
 sky130_fd_sc_hd__o211a_1 _8488_ (.A1(_3530_),
    .A2(_3601_),
    .B1(_3628_),
    .C1(_3350_),
    .X(_0074_));
 sky130_fd_sc_hd__o221a_1 _8489_ (.A1(_3315_),
    .A2(_3345_),
    .B1(_3621_),
    .B2(_3311_),
    .C1(_3534_),
    .X(_3629_));
 sky130_fd_sc_hd__o31a_1 _8490_ (.A1(_3307_),
    .A2(_3310_),
    .A3(_3589_),
    .B1(_3629_),
    .X(_3630_));
 sky130_fd_sc_hd__a221o_1 _8491_ (.A1(_3486_),
    .A2(_3418_),
    .B1(_3623_),
    .B2(_3311_),
    .C1(_3630_),
    .X(_3631_));
 sky130_fd_sc_hd__xor2_2 _8492_ (.A(net116),
    .B(_3631_),
    .X(_3632_));
 sky130_fd_sc_hd__nor2_1 _8493_ (.A(_3544_),
    .B(_3625_),
    .Y(_3633_));
 sky130_fd_sc_hd__a211o_1 _8494_ (.A1(_3544_),
    .A2(_3632_),
    .B1(_3633_),
    .C1(_3563_),
    .X(_3634_));
 sky130_fd_sc_hd__o211a_1 _8495_ (.A1(_3527_),
    .A2(_3617_),
    .B1(_3634_),
    .C1(_3350_),
    .X(_0075_));
 sky130_fd_sc_hd__nand2_1 _8496_ (.A(_3563_),
    .B(_3625_),
    .Y(_3636_));
 sky130_fd_sc_hd__a311o_1 _8497_ (.A1(_3330_),
    .A2(_3484_),
    .A3(_3618_),
    .B1(_3620_),
    .C1(_3329_),
    .X(_3637_));
 sky130_fd_sc_hd__mux2_1 _8498_ (.A0(_3318_),
    .A1(_3504_),
    .S(_3344_),
    .X(_3638_));
 sky130_fd_sc_hd__a21oi_1 _8499_ (.A1(_3416_),
    .A2(_3622_),
    .B1(_3421_),
    .Y(_3639_));
 sky130_fd_sc_hd__nor2_1 _8500_ (.A(_3569_),
    .B(_3639_),
    .Y(_3640_));
 sky130_fd_sc_hd__a31o_1 _8501_ (.A1(_3569_),
    .A2(_3637_),
    .A3(_3638_),
    .B1(_3640_),
    .X(_3641_));
 sky130_fd_sc_hd__xnor2_2 _8502_ (.A(net110),
    .B(_3641_),
    .Y(_3642_));
 sky130_fd_sc_hd__o21a_1 _8503_ (.A1(_3560_),
    .A2(_3642_),
    .B1(_3348_),
    .X(_3643_));
 sky130_fd_sc_hd__o211a_1 _8504_ (.A1(_3543_),
    .A2(_3632_),
    .B1(_3636_),
    .C1(_3643_),
    .X(_0076_));
 sky130_fd_sc_hd__inv_2 _8505_ (.A(_3320_),
    .Y(_3644_));
 sky130_fd_sc_hd__mux2_1 _8506_ (.A0(_3644_),
    .A1(_3508_),
    .S(_3589_),
    .X(_3646_));
 sky130_fd_sc_hd__a31o_1 _8507_ (.A1(_3287_),
    .A2(_3637_),
    .A3(_3638_),
    .B1(_3646_),
    .X(_3647_));
 sky130_fd_sc_hd__o21ai_1 _8508_ (.A1(_3287_),
    .A2(_3639_),
    .B1(_3424_),
    .Y(_3648_));
 sky130_fd_sc_hd__mux2_1 _8509_ (.A0(_3647_),
    .A1(_3648_),
    .S(_3486_),
    .X(_3649_));
 sky130_fd_sc_hd__xnor2_2 _8510_ (.A(_3649_),
    .B(_3293_),
    .Y(_3650_));
 sky130_fd_sc_hd__o221ai_1 _8511_ (.A1(_3530_),
    .A2(_3632_),
    .B1(_3560_),
    .B2(_3650_),
    .C1(_1676_),
    .Y(_3651_));
 sky130_fd_sc_hd__o21ba_1 _8512_ (.A1(_3543_),
    .A2(_3642_),
    .B1_N(_3651_),
    .X(_0077_));
 sky130_fd_sc_hd__o31ai_1 _8513_ (.A1(_3287_),
    .A2(_3293_),
    .A3(_3639_),
    .B1(_3428_),
    .Y(_3652_));
 sky130_fd_sc_hd__nand2_1 _8514_ (.A(_3287_),
    .B(_3293_),
    .Y(_3653_));
 sky130_fd_sc_hd__a21o_1 _8515_ (.A1(_3637_),
    .A2(_3638_),
    .B1(_3653_),
    .X(_3654_));
 sky130_fd_sc_hd__o211a_1 _8516_ (.A1(_3508_),
    .A2(_3322_),
    .B1(_3321_),
    .C1(_3344_),
    .X(_3656_));
 sky130_fd_sc_hd__a21oi_1 _8517_ (.A1(_3323_),
    .A2(_3589_),
    .B1(_3656_),
    .Y(_3657_));
 sky130_fd_sc_hd__and3_1 _8518_ (.A(_3535_),
    .B(_3654_),
    .C(_3657_),
    .X(_3658_));
 sky130_fd_sc_hd__a21o_1 _8519_ (.A1(_3486_),
    .A2(_3652_),
    .B1(_3658_),
    .X(_3659_));
 sky130_fd_sc_hd__xor2_2 _8520_ (.A(net129),
    .B(_3659_),
    .X(_3660_));
 sky130_fd_sc_hd__o22a_1 _8521_ (.A1(_3543_),
    .A2(_3650_),
    .B1(_3660_),
    .B2(_3560_),
    .X(_3661_));
 sky130_fd_sc_hd__o211a_1 _8522_ (.A1(_3530_),
    .A2(_3642_),
    .B1(_3661_),
    .C1(_3350_),
    .X(_0078_));
 sky130_fd_sc_hd__a21o_1 _8523_ (.A1(_3654_),
    .A2(_3657_),
    .B1(_3280_),
    .X(_3662_));
 sky130_fd_sc_hd__nand2_1 _8524_ (.A(_3276_),
    .B(_3279_),
    .Y(_3663_));
 sky130_fd_sc_hd__mux2_1 _8525_ (.A0(_3663_),
    .A1(_3506_),
    .S(_3345_),
    .X(_3664_));
 sky130_fd_sc_hd__a21oi_1 _8526_ (.A1(_3280_),
    .A2(_3652_),
    .B1(_3407_),
    .Y(_3666_));
 sky130_fd_sc_hd__nor2_1 _8527_ (.A(_3569_),
    .B(_3666_),
    .Y(_3667_));
 sky130_fd_sc_hd__a31o_1 _8528_ (.A1(_3569_),
    .A2(_3662_),
    .A3(_3664_),
    .B1(_3667_),
    .X(_3668_));
 sky130_fd_sc_hd__xnor2_2 _8529_ (.A(_3273_),
    .B(_3668_),
    .Y(_3669_));
 sky130_fd_sc_hd__o221a_1 _8530_ (.A1(_3529_),
    .A2(_3650_),
    .B1(_3660_),
    .B2(_3543_),
    .C1(_3348_),
    .X(_3670_));
 sky130_fd_sc_hd__a21boi_1 _8531_ (.A1(_3544_),
    .A2(_3669_),
    .B1_N(_3670_),
    .Y(_0079_));
 sky130_fd_sc_hd__nand2_1 _8532_ (.A(_3431_),
    .B(_3463_),
    .Y(_3671_));
 sky130_fd_sc_hd__o211a_1 _8533_ (.A1(_2818_),
    .A2(_3339_),
    .B1(_3511_),
    .C1(_3343_),
    .X(_3672_));
 sky130_fd_sc_hd__a21oi_1 _8534_ (.A1(_3333_),
    .A2(_3484_),
    .B1(_3672_),
    .Y(_3673_));
 sky130_fd_sc_hd__mux2_1 _8535_ (.A0(_3671_),
    .A1(_3673_),
    .S(_3534_),
    .X(_3674_));
 sky130_fd_sc_hd__xnor2_2 _8536_ (.A(_2932_),
    .B(_3674_),
    .Y(_3676_));
 sky130_fd_sc_hd__inv_2 _8537_ (.A(_3676_),
    .Y(_3677_));
 sky130_fd_sc_hd__nand2_1 _8538_ (.A(_3553_),
    .B(_3669_),
    .Y(_3678_));
 sky130_fd_sc_hd__or2_1 _8539_ (.A(net133),
    .B(_3660_),
    .X(_3679_));
 sky130_fd_sc_hd__o2111a_1 _8540_ (.A1(_3560_),
    .A2(_3677_),
    .B1(_3678_),
    .C1(_1676_),
    .D1(_3679_),
    .X(_0080_));
 sky130_fd_sc_hd__o221a_1 _8541_ (.A1(_2929_),
    .A2(_3345_),
    .B1(_3673_),
    .B2(_2932_),
    .C1(_3534_),
    .X(_3680_));
 sky130_fd_sc_hd__o21a_1 _8542_ (.A1(_2930_),
    .A2(_3589_),
    .B1(_3680_),
    .X(_3681_));
 sky130_fd_sc_hd__nand2_1 _8543_ (.A(_2932_),
    .B(_3671_),
    .Y(_3682_));
 sky130_fd_sc_hd__a21oi_1 _8544_ (.A1(_3682_),
    .A2(_3468_),
    .B1(_3569_),
    .Y(_3683_));
 sky130_fd_sc_hd__nor2_1 _8545_ (.A(_3681_),
    .B(_3683_),
    .Y(_3684_));
 sky130_fd_sc_hd__xnor2_2 _8546_ (.A(_2904_),
    .B(_3684_),
    .Y(_3686_));
 sky130_fd_sc_hd__o221a_1 _8547_ (.A1(_3524_),
    .A2(_3677_),
    .B1(_3686_),
    .B2(_3560_),
    .C1(_3348_),
    .X(_3687_));
 sky130_fd_sc_hd__a21boi_1 _8548_ (.A1(_3563_),
    .A2(_3669_),
    .B1_N(_3687_),
    .Y(_0081_));
 sky130_fd_sc_hd__nand2_1 _8549_ (.A(_3563_),
    .B(_3676_),
    .Y(_3688_));
 sky130_fd_sc_hd__o21ai_1 _8550_ (.A1(_3464_),
    .A2(_3682_),
    .B1(_3471_),
    .Y(_3689_));
 sky130_fd_sc_hd__inv_2 _8551_ (.A(_2933_),
    .Y(_3690_));
 sky130_fd_sc_hd__nand2_1 _8552_ (.A(_3336_),
    .B(_3589_),
    .Y(_3691_));
 sky130_fd_sc_hd__o221a_1 _8553_ (.A1(_3589_),
    .A2(_3513_),
    .B1(_3673_),
    .B2(_3690_),
    .C1(_3691_),
    .X(_3692_));
 sky130_fd_sc_hd__mux2_1 _8554_ (.A0(_3689_),
    .A1(_3692_),
    .S(_3569_),
    .X(_3693_));
 sky130_fd_sc_hd__xnor2_2 _8555_ (.A(_2877_),
    .B(_3693_),
    .Y(_3694_));
 sky130_fd_sc_hd__nand2_1 _8556_ (.A(_3544_),
    .B(_3694_),
    .Y(_3696_));
 sky130_fd_sc_hd__o2111a_1 _8557_ (.A1(_3543_),
    .A2(_3686_),
    .B1(_3688_),
    .C1(_3696_),
    .D1(_1676_),
    .X(_0082_));
 sky130_fd_sc_hd__a21o_1 _8558_ (.A1(_2877_),
    .A2(_3689_),
    .B1(_3473_),
    .X(_3697_));
 sky130_fd_sc_hd__mux2_1 _8559_ (.A0(_2874_),
    .A1(_2875_),
    .S(_3345_),
    .X(_3698_));
 sky130_fd_sc_hd__o211a_1 _8560_ (.A1(_2877_),
    .A2(_3692_),
    .B1(_3698_),
    .C1(_3535_),
    .X(_3699_));
 sky130_fd_sc_hd__a21oi_1 _8561_ (.A1(_3486_),
    .A2(_3697_),
    .B1(_3699_),
    .Y(_3700_));
 sky130_fd_sc_hd__xnor2_2 _8562_ (.A(_2848_),
    .B(_3700_),
    .Y(_3701_));
 sky130_fd_sc_hd__o221a_1 _8563_ (.A1(net133),
    .A2(_3686_),
    .B1(_3701_),
    .B2(_3560_),
    .C1(_3348_),
    .X(_3702_));
 sky130_fd_sc_hd__a21boi_1 _8564_ (.A1(_3553_),
    .A2(_3694_),
    .B1_N(_3702_),
    .Y(_0083_));
 sky130_fd_sc_hd__nand2_1 _8565_ (.A(_3467_),
    .B(_3476_),
    .Y(_3703_));
 sky130_fd_sc_hd__a21oi_1 _8566_ (.A1(net103),
    .A2(_3589_),
    .B1(_3518_),
    .Y(_3705_));
 sky130_fd_sc_hd__nand2_1 _8567_ (.A(_3569_),
    .B(_3705_),
    .Y(_3706_));
 sky130_fd_sc_hd__o21a_1 _8568_ (.A1(_3569_),
    .A2(_3703_),
    .B1(_3706_),
    .X(_3707_));
 sky130_fd_sc_hd__xnor2_2 _8569_ (.A(_3479_),
    .B(_3707_),
    .Y(_3708_));
 sky130_fd_sc_hd__o221a_1 _8570_ (.A1(_3524_),
    .A2(_3701_),
    .B1(_3708_),
    .B2(_3559_),
    .C1(_3348_),
    .X(_3709_));
 sky130_fd_sc_hd__a21boi_1 _8571_ (.A1(_3563_),
    .A2(_3694_),
    .B1_N(_3709_),
    .Y(_0084_));
 sky130_fd_sc_hd__mux2_1 _8572_ (.A0(_2791_),
    .A1(_2792_),
    .S(_3589_),
    .X(_3710_));
 sky130_fd_sc_hd__o21ai_1 _8573_ (.A1(_2793_),
    .A2(_3705_),
    .B1(_3710_),
    .Y(_3711_));
 sky130_fd_sc_hd__a211o_1 _8574_ (.A1(_2793_),
    .A2(_3703_),
    .B1(_3395_),
    .C1(_3534_),
    .X(_3712_));
 sky130_fd_sc_hd__o21a_1 _8575_ (.A1(_3486_),
    .A2(_3711_),
    .B1(_3712_),
    .X(_3713_));
 sky130_fd_sc_hd__xnor2_1 _8576_ (.A(_2816_),
    .B(_3713_),
    .Y(_3715_));
 sky130_fd_sc_hd__nand2_1 _8577_ (.A(_3544_),
    .B(_3715_),
    .Y(_3716_));
 sky130_fd_sc_hd__o21a_1 _8578_ (.A1(_3530_),
    .A2(_3701_),
    .B1(_3348_),
    .X(_3717_));
 sky130_fd_sc_hd__o211a_1 _8579_ (.A1(_3543_),
    .A2(_3708_),
    .B1(_3716_),
    .C1(_3717_),
    .X(_0085_));
 sky130_fd_sc_hd__a311o_1 _8580_ (.A1(_2793_),
    .A2(_2816_),
    .A3(_3703_),
    .B1(_3398_),
    .C1(_3535_),
    .X(_3718_));
 sky130_fd_sc_hd__and3_1 _8581_ (.A(_3490_),
    .B(_3519_),
    .C(_3718_),
    .X(_3719_));
 sky130_fd_sc_hd__xnor2_1 _8582_ (.A(_2752_),
    .B(_3719_),
    .Y(_3720_));
 sky130_fd_sc_hd__nor2_1 _8583_ (.A(net111),
    .B(_3715_),
    .Y(_3721_));
 sky130_fd_sc_hd__a211o_1 _8584_ (.A1(_3544_),
    .A2(_3720_),
    .B1(_3721_),
    .C1(_3563_),
    .X(_3722_));
 sky130_fd_sc_hd__o211a_1 _8585_ (.A1(_3530_),
    .A2(_3708_),
    .B1(_3722_),
    .C1(_3350_),
    .X(_0086_));
 sky130_fd_sc_hd__o221a_1 _8586_ (.A1(_3527_),
    .A2(_3721_),
    .B1(_3720_),
    .B2(_3543_),
    .C1(_3350_),
    .X(_0087_));
 sky130_fd_sc_hd__or2_2 _8587_ (.A(_2697_),
    .B(_2698_),
    .X(_3724_));
 sky130_fd_sc_hd__or3_1 _8588_ (.A(_3724_),
    .B(net111),
    .C(_3527_),
    .X(_3725_));
 sky130_fd_sc_hd__xnor2_1 _8589_ (.A(_3724_),
    .B(_3559_),
    .Y(_3726_));
 sky130_fd_sc_hd__nand2_1 _8590_ (.A(_3530_),
    .B(_3726_),
    .Y(_3727_));
 sky130_fd_sc_hd__a21oi_1 _8591_ (.A1(_3725_),
    .A2(_3727_),
    .B1(_3597_),
    .Y(_0088_));
 sky130_fd_sc_hd__nor2_1 _8592_ (.A(_2635_),
    .B(_2831_),
    .Y(_3728_));
 sky130_fd_sc_hd__a31o_1 _8593_ (.A1(_2627_),
    .A2(_2636_),
    .A3(_2831_),
    .B1(_3728_),
    .X(_3729_));
 sky130_fd_sc_hd__nand2_1 _8594_ (.A(_3724_),
    .B(_3729_),
    .Y(_3730_));
 sky130_fd_sc_hd__or2_1 _8595_ (.A(_3724_),
    .B(_3729_),
    .X(_3731_));
 sky130_fd_sc_hd__and2_1 _8596_ (.A(_3730_),
    .B(_3731_),
    .X(_3733_));
 sky130_fd_sc_hd__mux2_4 _8597_ (.A0(_3729_),
    .A1(_3733_),
    .S(_3482_),
    .X(_3734_));
 sky130_fd_sc_hd__or3_4 _8598_ (.A(net111),
    .B(_3527_),
    .C(_3731_),
    .X(_3735_));
 sky130_fd_sc_hd__a21bo_1 _8599_ (.A1(_3725_),
    .A2(_3734_),
    .B1_N(_3735_),
    .X(_3736_));
 sky130_fd_sc_hd__and2_1 _8600_ (.A(_3383_),
    .B(_3736_),
    .X(_3737_));
 sky130_fd_sc_hd__clkbuf_1 _8601_ (.A(_3737_),
    .X(_0089_));
 sky130_fd_sc_hd__a211o_1 _8602_ (.A1(_3405_),
    .A2(_3480_),
    .B1(_3730_),
    .C1(_3534_),
    .X(_3738_));
 sky130_fd_sc_hd__mux2_1 _8603_ (.A0(_2628_),
    .A1(net83),
    .S(_2748_),
    .X(_3739_));
 sky130_fd_sc_hd__xnor2_1 _8604_ (.A(_3738_),
    .B(_3739_),
    .Y(_3740_));
 sky130_fd_sc_hd__or3_1 _8605_ (.A(_3726_),
    .B(_3734_),
    .C(_3740_),
    .X(_3741_));
 sky130_fd_sc_hd__a2bb2o_1 _8606_ (.A1_N(_3529_),
    .A2_N(_3741_),
    .B1(_3740_),
    .B2(_3735_),
    .X(_3743_));
 sky130_fd_sc_hd__and2_1 _8607_ (.A(_3383_),
    .B(_3743_),
    .X(_3744_));
 sky130_fd_sc_hd__clkbuf_1 _8608_ (.A(_3744_),
    .X(_0090_));
 sky130_fd_sc_hd__inv_2 _8609_ (.A(_2621_),
    .Y(_3745_));
 sky130_fd_sc_hd__mux2_1 _8610_ (.A0(_3745_),
    .A1(net84),
    .S(_2748_),
    .X(_3746_));
 sky130_fd_sc_hd__and2_1 _8611_ (.A(_3739_),
    .B(_3746_),
    .X(_3747_));
 sky130_fd_sc_hd__nand2b_1 _8612_ (.A_N(_3738_),
    .B(_3747_),
    .Y(_3748_));
 sky130_fd_sc_hd__and2_1 _8613_ (.A(_3724_),
    .B(_3729_),
    .X(_3749_));
 sky130_fd_sc_hd__a31o_1 _8614_ (.A1(_3482_),
    .A2(_3749_),
    .A3(_3739_),
    .B1(_3746_),
    .X(_3750_));
 sky130_fd_sc_hd__o211a_1 _8615_ (.A1(net133),
    .A2(_3741_),
    .B1(_3748_),
    .C1(_3750_),
    .X(_3751_));
 sky130_fd_sc_hd__a2111oi_4 _8616_ (.A1(_3748_),
    .A2(_3750_),
    .B1(_3726_),
    .C1(_3734_),
    .D1(_3740_),
    .Y(_3753_));
 sky130_fd_sc_hd__and2_4 _8617_ (.A(_3562_),
    .B(_3753_),
    .X(_3754_));
 sky130_fd_sc_hd__o21a_1 _8618_ (.A1(_3751_),
    .A2(_3754_),
    .B1(_3350_),
    .X(_0091_));
 sky130_fd_sc_hd__nor2_1 _8619_ (.A(_2600_),
    .B(_2748_),
    .Y(_3755_));
 sky130_fd_sc_hd__a21o_1 _8620_ (.A1(net85),
    .A2(_2748_),
    .B1(_3755_),
    .X(_3756_));
 sky130_fd_sc_hd__a31oi_1 _8621_ (.A1(_3482_),
    .A2(_3749_),
    .A3(_3747_),
    .B1(_3756_),
    .Y(_3757_));
 sky130_fd_sc_hd__nand2_1 _8622_ (.A(_3747_),
    .B(_3756_),
    .Y(_3758_));
 sky130_fd_sc_hd__nor2_1 _8623_ (.A(_3738_),
    .B(_3758_),
    .Y(_3759_));
 sky130_fd_sc_hd__or2_1 _8624_ (.A(_3757_),
    .B(_3759_),
    .X(_3760_));
 sky130_fd_sc_hd__xor2_1 _8625_ (.A(_3754_),
    .B(_3760_),
    .X(_3761_));
 sky130_fd_sc_hd__nor2_1 _8626_ (.A(_3597_),
    .B(_3761_),
    .Y(_0092_));
 sky130_fd_sc_hd__a2111o_1 _8627_ (.A1(_3405_),
    .A2(_3480_),
    .B1(_3730_),
    .C1(_3758_),
    .D1(_3534_),
    .X(_3763_));
 sky130_fd_sc_hd__and3_1 _8628_ (.A(_2585_),
    .B(_2597_),
    .C(_2831_),
    .X(_3764_));
 sky130_fd_sc_hd__a21o_1 _8629_ (.A1(net86),
    .A2(_2748_),
    .B1(_3764_),
    .X(_3765_));
 sky130_fd_sc_hd__xor2_1 _8630_ (.A(_3763_),
    .B(_3765_),
    .X(_3766_));
 sky130_fd_sc_hd__a21oi_1 _8631_ (.A1(_3754_),
    .A2(_3760_),
    .B1(_3766_),
    .Y(_3767_));
 sky130_fd_sc_hd__and4_1 _8632_ (.A(_3753_),
    .B(_3562_),
    .C(_3760_),
    .D(_3766_),
    .X(_3768_));
 sky130_fd_sc_hd__o21a_1 _8633_ (.A1(_3767_),
    .A2(_3768_),
    .B1(_3350_),
    .X(_0093_));
 sky130_fd_sc_hd__nand2b_1 _8634_ (.A_N(_3763_),
    .B(_3765_),
    .Y(_3769_));
 sky130_fd_sc_hd__inv_2 _8635_ (.A(net87),
    .Y(_3770_));
 sky130_fd_sc_hd__mux2_1 _8636_ (.A0(_2592_),
    .A1(_3770_),
    .S(_2748_),
    .X(_3772_));
 sky130_fd_sc_hd__xor2_1 _8637_ (.A(_3769_),
    .B(_3772_),
    .X(_3773_));
 sky130_fd_sc_hd__xnor2_1 _8638_ (.A(_3768_),
    .B(_3773_),
    .Y(_3774_));
 sky130_fd_sc_hd__nor2_1 _8639_ (.A(_3597_),
    .B(_3774_),
    .Y(_0094_));
 sky130_fd_sc_hd__o21ai_1 _8640_ (.A1(_3757_),
    .A2(_3759_),
    .B1(_3766_),
    .Y(_3775_));
 sky130_fd_sc_hd__and4bb_1 _8641_ (.A_N(_3773_),
    .B_N(_3775_),
    .C(_3753_),
    .D(_3562_),
    .X(_3776_));
 sky130_fd_sc_hd__or2_1 _8642_ (.A(_3769_),
    .B(_3772_),
    .X(_3777_));
 sky130_fd_sc_hd__nor2_1 _8643_ (.A(_2607_),
    .B(net114),
    .Y(_3778_));
 sky130_fd_sc_hd__a31o_1 _8644_ (.A1(_3778_),
    .A2(_2654_),
    .A3(_2695_),
    .B1(net89),
    .X(_3779_));
 sky130_fd_sc_hd__xnor2_1 _8645_ (.A(_3777_),
    .B(_3779_),
    .Y(_3780_));
 sky130_fd_sc_hd__xnor2_1 _8646_ (.A(_3776_),
    .B(_3780_),
    .Y(_3782_));
 sky130_fd_sc_hd__nor2_1 _8647_ (.A(_3597_),
    .B(_3782_),
    .Y(_0095_));
 sky130_fd_sc_hd__dfxtp_1 _8648_ (.CLK(clknet_3_5__leaf_CLK),
    .D(_0000_),
    .Q(\In1_reg[0] ));
 sky130_fd_sc_hd__dfxtp_4 _8649_ (.CLK(clknet_3_5__leaf_CLK),
    .D(_0001_),
    .Q(\In1_reg[1] ));
 sky130_fd_sc_hd__dfxtp_2 _8650_ (.CLK(clknet_3_5__leaf_CLK),
    .D(_0002_),
    .Q(\In1_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _8651_ (.CLK(clknet_3_5__leaf_CLK),
    .D(_0003_),
    .Q(\In1_reg[3] ));
 sky130_fd_sc_hd__dfxtp_4 _8652_ (.CLK(clknet_3_3__leaf_CLK),
    .D(_0004_),
    .Q(\In1_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8653_ (.CLK(clknet_3_5__leaf_CLK),
    .D(_0005_),
    .Q(\In1_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8654_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0006_),
    .Q(\In1_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8655_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0007_),
    .Q(\In1_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8656_ (.CLK(clknet_3_4__leaf_CLK),
    .D(_0008_),
    .Q(\In1_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8657_ (.CLK(clknet_3_4__leaf_CLK),
    .D(_0009_),
    .Q(\In1_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8658_ (.CLK(clknet_3_4__leaf_CLK),
    .D(_0010_),
    .Q(\In1_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8659_ (.CLK(clknet_3_4__leaf_CLK),
    .D(_0011_),
    .Q(\In1_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8660_ (.CLK(clknet_3_4__leaf_CLK),
    .D(_0012_),
    .Q(\In1_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8661_ (.CLK(clknet_3_4__leaf_CLK),
    .D(_0013_),
    .Q(\In1_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8662_ (.CLK(clknet_3_3__leaf_CLK),
    .D(_0014_),
    .Q(\In1_reg[14] ));
 sky130_fd_sc_hd__dfxtp_2 _8663_ (.CLK(clknet_3_3__leaf_CLK),
    .D(_0015_),
    .Q(\In1_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8664_ (.CLK(clknet_3_4__leaf_CLK),
    .D(_0016_),
    .Q(\In1_reg[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8665_ (.CLK(clknet_3_4__leaf_CLK),
    .D(_0017_),
    .Q(\In1_reg[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8666_ (.CLK(clknet_3_3__leaf_CLK),
    .D(_0018_),
    .Q(\In1_reg[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8667_ (.CLK(clknet_3_4__leaf_CLK),
    .D(_0019_),
    .Q(\In1_reg[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8668_ (.CLK(clknet_3_0__leaf_CLK),
    .D(_0020_),
    .Q(\In1_reg[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8669_ (.CLK(clknet_3_4__leaf_CLK),
    .D(_0021_),
    .Q(\In1_reg[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8670_ (.CLK(clknet_3_0__leaf_CLK),
    .D(_0022_),
    .Q(\In1_reg[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8671_ (.CLK(clknet_3_3__leaf_CLK),
    .D(_0023_),
    .Q(\M1.ua1.fa0.a ));
 sky130_fd_sc_hd__dfxtp_1 _8672_ (.CLK(clknet_3_3__leaf_CLK),
    .D(_0024_),
    .Q(\M1.ua1.fa1.a ));
 sky130_fd_sc_hd__dfxtp_1 _8673_ (.CLK(clknet_3_3__leaf_CLK),
    .D(_0025_),
    .Q(\M1.ua1.fa2.a ));
 sky130_fd_sc_hd__dfxtp_1 _8674_ (.CLK(clknet_3_3__leaf_CLK),
    .D(_0026_),
    .Q(\M1.ua1.fa3.a ));
 sky130_fd_sc_hd__dfxtp_1 _8675_ (.CLK(clknet_3_3__leaf_CLK),
    .D(_0027_),
    .Q(\M1.ua1.fa4.a ));
 sky130_fd_sc_hd__dfxtp_1 _8676_ (.CLK(clknet_3_3__leaf_CLK),
    .D(_0028_),
    .Q(\M1.ua1.fa5.a ));
 sky130_fd_sc_hd__dfxtp_1 _8677_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0029_),
    .Q(\M1.ua1.fa6.a ));
 sky130_fd_sc_hd__dfxtp_1 _8678_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0030_),
    .Q(\M1.ua1.fa7.a ));
 sky130_fd_sc_hd__dfxtp_1 _8679_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0031_),
    .Q(\In1_reg[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8680_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0032_),
    .Q(\F1.sign_b ));
 sky130_fd_sc_hd__dfxtp_2 _8681_ (.CLK(clknet_3_5__leaf_CLK),
    .D(_0033_),
    .Q(\In2_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8682_ (.CLK(clknet_3_5__leaf_CLK),
    .D(_0034_),
    .Q(\M1.U1.U1.u2.instance9_8.Prop_L ));
 sky130_fd_sc_hd__dfxtp_2 _8683_ (.CLK(clknet_3_5__leaf_CLK),
    .D(_0035_),
    .Q(\In2_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8684_ (.CLK(clknet_3_5__leaf_CLK),
    .D(_0036_),
    .Q(\M1.U1.U2.u2.instance11_10.Prop_L ));
 sky130_fd_sc_hd__dfxtp_1 _8685_ (.CLK(clknet_3_6__leaf_CLK),
    .D(_0037_),
    .Q(\In2_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8686_ (.CLK(clknet_3_6__leaf_CLK),
    .D(_0038_),
    .Q(\M1.U1.U3.u2.instance13_12.Prop_L ));
 sky130_fd_sc_hd__dfxtp_1 _8687_ (.CLK(clknet_3_6__leaf_CLK),
    .D(_0039_),
    .Q(\In2_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8688_ (.CLK(clknet_3_6__leaf_CLK),
    .D(_0040_),
    .Q(\M1.U1.U4.u2.instance15_14.Prop_L ));
 sky130_fd_sc_hd__dfxtp_1 _8689_ (.CLK(clknet_3_7__leaf_CLK),
    .D(_0041_),
    .Q(\In2_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8690_ (.CLK(clknet_3_6__leaf_CLK),
    .D(_0042_),
    .Q(\M1.U1.U5.u3.instance1_0.Prop_L ));
 sky130_fd_sc_hd__dfxtp_1 _8691_ (.CLK(clknet_3_7__leaf_CLK),
    .D(_0043_),
    .Q(\In2_reg[10] ));
 sky130_fd_sc_hd__dfxtp_2 _8692_ (.CLK(clknet_3_7__leaf_CLK),
    .D(_0044_),
    .Q(\M1.U1.U6.u3.instance3_2.Prop_L ));
 sky130_fd_sc_hd__dfxtp_1 _8693_ (.CLK(clknet_3_7__leaf_CLK),
    .D(_0045_),
    .Q(\In2_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8694_ (.CLK(clknet_3_7__leaf_CLK),
    .D(_0046_),
    .Q(\M1.U1.U7.u3.instance5_4.Prop_L ));
 sky130_fd_sc_hd__dfxtp_1 _8695_ (.CLK(clknet_3_7__leaf_CLK),
    .D(_0047_),
    .Q(\In2_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8696_ (.CLK(clknet_3_7__leaf_CLK),
    .D(_0048_),
    .Q(\M1.U1.U8.u3.instance7_6.Prop_L ));
 sky130_fd_sc_hd__dfxtp_1 _8697_ (.CLK(clknet_3_7__leaf_CLK),
    .D(_0049_),
    .Q(\In2_reg[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8698_ (.CLK(clknet_3_6__leaf_CLK),
    .D(_0050_),
    .Q(\M1.U1.U9.u3.instance9_8.Prop_L ));
 sky130_fd_sc_hd__dfxtp_1 _8699_ (.CLK(clknet_3_6__leaf_CLK),
    .D(_0051_),
    .Q(\In2_reg[18] ));
 sky130_fd_sc_hd__dfxtp_2 _8700_ (.CLK(clknet_3_7__leaf_CLK),
    .D(_0052_),
    .Q(\M1.U1.U10.u3.instance11_10.Prop_L ));
 sky130_fd_sc_hd__dfxtp_1 _8701_ (.CLK(clknet_3_6__leaf_CLK),
    .D(_0053_),
    .Q(\In2_reg[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8702_ (.CLK(clknet_3_7__leaf_CLK),
    .D(_0054_),
    .Q(\M1.U1.U11.u3.instance13_12.Prop_L ));
 sky130_fd_sc_hd__dfxtp_2 _8703_ (.CLK(clknet_3_7__leaf_CLK),
    .D(_0055_),
    .Q(\In2_reg[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8704_ (.CLK(clknet_3_5__leaf_CLK),
    .D(_0056_),
    .Q(\M1.ua1.fa0.b ));
 sky130_fd_sc_hd__dfxtp_1 _8705_ (.CLK(clknet_3_3__leaf_CLK),
    .D(_0057_),
    .Q(\M1.ua1.fa1.b ));
 sky130_fd_sc_hd__dfxtp_1 _8706_ (.CLK(clknet_3_3__leaf_CLK),
    .D(_0058_),
    .Q(\M1.ua1.fa2.b ));
 sky130_fd_sc_hd__dfxtp_1 _8707_ (.CLK(clknet_3_3__leaf_CLK),
    .D(_0059_),
    .Q(\M1.ua1.fa3.b ));
 sky130_fd_sc_hd__dfxtp_1 _8708_ (.CLK(clknet_3_3__leaf_CLK),
    .D(_0060_),
    .Q(\M1.ua1.fa4.b ));
 sky130_fd_sc_hd__dfxtp_1 _8709_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0061_),
    .Q(\M1.ua1.fa5.b ));
 sky130_fd_sc_hd__dfxtp_1 _8710_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0062_),
    .Q(\M1.ua1.fa6.b ));
 sky130_fd_sc_hd__dfxtp_1 _8711_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0063_),
    .Q(\M1.ua1.fa7.b ));
 sky130_fd_sc_hd__dfxtp_1 _8712_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0064_),
    .Q(\In2_reg[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8713_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_0065_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_1 _8714_ (.CLK(clknet_3_0__leaf_CLK),
    .D(_0066_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_2 _8715_ (.CLK(clknet_3_0__leaf_CLK),
    .D(_0067_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_2 _8716_ (.CLK(clknet_3_0__leaf_CLK),
    .D(_0068_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_2 _8717_ (.CLK(clknet_3_0__leaf_CLK),
    .D(_0069_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_2 _8718_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_0070_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_2 _8719_ (.CLK(clknet_3_0__leaf_CLK),
    .D(_0071_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_2 _8720_ (.CLK(clknet_3_0__leaf_CLK),
    .D(_0072_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_1 _8721_ (.CLK(clknet_3_0__leaf_CLK),
    .D(_0073_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _8722_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_0074_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_1 _8723_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_0075_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _8724_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_0076_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_2 _8725_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_0077_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_1 _8726_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_0078_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_1 _8727_ (.CLK(clknet_3_0__leaf_CLK),
    .D(_0079_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_1 _8728_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_0080_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_1 _8729_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_0081_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _8730_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_0082_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _8731_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_0083_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_2 _8732_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_0084_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_1 _8733_ (.CLK(clknet_3_1__leaf_CLK),
    .D(_0085_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_2 _8734_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0086_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_1 _8735_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0087_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_4 _8736_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0088_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_1 _8737_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0089_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_2 _8738_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0090_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_1 _8739_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0091_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_2 _8740_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0092_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_1 _8741_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0093_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_1 _8742_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0094_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_2 _8743_ (.CLK(clknet_3_2__leaf_CLK),
    .D(_0095_),
    .Q(net89));
 sky130_fd_sc_hd__clkbuf_1 _8744_ (.A(\F1.sign_b ),
    .X(net90));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1507 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(In1[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(In1[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(In1[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(In1[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(In1[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(In1[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(In1[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(In1[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(In1[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(In1[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(In1[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(In1[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(In1[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(In1[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(In1[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(In1[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(In1[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(In1[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(In1[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(In1[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(In1[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(In1[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(In1[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(In1[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(In1[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(In1[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(In1[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(In1[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(In1[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(In1[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(In1[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(In1[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(In2[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(In2[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(In2[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(In2[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(In2[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(In2[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(In2[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(In2[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(In2[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(In2[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(In2[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(In2[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(In2[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(In2[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(In2[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(In2[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(In2[24]),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 input50 (.A(In2[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(In2[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(In2[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(In2[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(In2[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(In2[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(In2[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(In2[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(In2[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(In2[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(In2[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(In2[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(In2[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(In2[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(In2[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_8 input65 (.A(rst),
    .X(net65));
 sky130_fd_sc_hd__buf_1 output66 (.A(net66),
    .X(MacOut[0]));
 sky130_fd_sc_hd__buf_1 output67 (.A(net67),
    .X(MacOut[10]));
 sky130_fd_sc_hd__buf_1 output68 (.A(net68),
    .X(MacOut[11]));
 sky130_fd_sc_hd__buf_1 output69 (.A(net69),
    .X(MacOut[12]));
 sky130_fd_sc_hd__buf_1 output70 (.A(net70),
    .X(MacOut[13]));
 sky130_fd_sc_hd__buf_1 output71 (.A(net71),
    .X(MacOut[14]));
 sky130_fd_sc_hd__buf_1 output72 (.A(net72),
    .X(MacOut[15]));
 sky130_fd_sc_hd__buf_1 output73 (.A(net73),
    .X(MacOut[16]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net74),
    .X(MacOut[17]));
 sky130_fd_sc_hd__buf_1 output75 (.A(net75),
    .X(MacOut[18]));
 sky130_fd_sc_hd__buf_1 output76 (.A(net76),
    .X(MacOut[19]));
 sky130_fd_sc_hd__buf_1 output77 (.A(net77),
    .X(MacOut[1]));
 sky130_fd_sc_hd__buf_1 output78 (.A(net78),
    .X(MacOut[20]));
 sky130_fd_sc_hd__buf_1 output79 (.A(net79),
    .X(MacOut[21]));
 sky130_fd_sc_hd__buf_1 output80 (.A(net80),
    .X(MacOut[22]));
 sky130_fd_sc_hd__buf_1 output81 (.A(net81),
    .X(MacOut[23]));
 sky130_fd_sc_hd__buf_1 output82 (.A(net82),
    .X(MacOut[24]));
 sky130_fd_sc_hd__buf_1 output83 (.A(net83),
    .X(MacOut[25]));
 sky130_fd_sc_hd__buf_1 output84 (.A(net84),
    .X(MacOut[26]));
 sky130_fd_sc_hd__buf_1 output85 (.A(net85),
    .X(MacOut[27]));
 sky130_fd_sc_hd__buf_1 output86 (.A(net86),
    .X(MacOut[28]));
 sky130_fd_sc_hd__buf_1 output87 (.A(net87),
    .X(MacOut[29]));
 sky130_fd_sc_hd__buf_1 output88 (.A(net88),
    .X(MacOut[2]));
 sky130_fd_sc_hd__buf_1 output89 (.A(net89),
    .X(MacOut[30]));
 sky130_fd_sc_hd__buf_1 output90 (.A(net90),
    .X(MacOut[31]));
 sky130_fd_sc_hd__buf_1 output91 (.A(net91),
    .X(MacOut[3]));
 sky130_fd_sc_hd__buf_1 output92 (.A(net92),
    .X(MacOut[4]));
 sky130_fd_sc_hd__buf_1 output93 (.A(net93),
    .X(MacOut[5]));
 sky130_fd_sc_hd__buf_1 output94 (.A(net94),
    .X(MacOut[6]));
 sky130_fd_sc_hd__buf_1 output95 (.A(net95),
    .X(MacOut[7]));
 sky130_fd_sc_hd__buf_1 output96 (.A(net96),
    .X(MacOut[8]));
 sky130_fd_sc_hd__buf_1 output97 (.A(net97),
    .X(MacOut[9]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_CLK (.A(CLK),
    .X(clknet_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_0__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_1__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_2__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_3__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_4__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_5__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_6__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_7__leaf_CLK));
 sky130_fd_sc_hd__inv_8 clkload0 (.A(clknet_3_0__leaf_CLK));
 sky130_fd_sc_hd__clkinv_4 clkload1 (.A(clknet_3_1__leaf_CLK));
 sky130_fd_sc_hd__clkinv_4 clkload2 (.A(clknet_3_3__leaf_CLK));
 sky130_fd_sc_hd__inv_8 clkload3 (.A(clknet_3_4__leaf_CLK));
 sky130_fd_sc_hd__inv_8 clkload4 (.A(clknet_3_5__leaf_CLK));
 sky130_fd_sc_hd__clkinv_8 clkload5 (.A(clknet_3_6__leaf_CLK));
 sky130_fd_sc_hd__inv_6 clkload6 (.A(clknet_3_7__leaf_CLK));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(_2691_),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(_2691_),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(_2692_),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(_2602_),
    .X(net101));
 sky130_fd_sc_hd__buf_6 rebuffer5 (.A(_3339_),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net102),
    .X(net103));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer7 (.A(net102),
    .X(net104));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer8 (.A(_2317_),
    .X(net105));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer9 (.A(_2714_),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(_2639_),
    .X(net107));
 sky130_fd_sc_hd__buf_2 rebuffer11 (.A(_2640_),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(_2699_),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(_3287_),
    .X(net110));
 sky130_fd_sc_hd__a21oi_2 clone14 (.A1(_3480_),
    .A2(_3405_),
    .B1(_3401_),
    .Y(net111));
 sky130_fd_sc_hd__clkbuf_1 rebuffer15 (.A(_3165_),
    .X(net112));
 sky130_fd_sc_hd__buf_2 clone16 (.A(net115),
    .X(net113));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer17 (.A(_2615_),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(_2699_),
    .X(net115));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer19 (.A(_3303_),
    .X(net116));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer20 (.A(_2695_),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(_2695_),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(_2642_),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net119),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net119),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net125),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(_2760_),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer28 (.A(_2760_),
    .X(net125));
 sky130_fd_sc_hd__buf_4 split29 (.A(\In1_reg[1] ),
    .X(net126));
 sky130_fd_sc_hd__buf_2 rebuffer30 (.A(_2637_),
    .X(net127));
 sky130_fd_sc_hd__buf_6 rebuffer31 (.A(_2553_),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(_3280_),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(_2663_),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(_2663_),
    .X(net131));
 sky130_fd_sc_hd__buf_2 clone35 (.A(_2714_),
    .X(net132));
 sky130_fd_sc_hd__buf_2 clone36 (.A(_3528_),
    .X(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_3171_));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_649 ();
endmodule
